//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_;
  NOR2_X1   g000(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NOR3_X1   g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT9), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(KEYINPUT9), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT10), .B(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n213_), .A2(new_n215_), .A3(G99gat), .A4(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n207_), .A2(new_n211_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n210_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n222_), .A2(new_n226_), .A3(new_n223_), .A4(new_n210_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n220_), .A2(new_n216_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n206_), .A2(KEYINPUT67), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n221_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G57gat), .B(G64gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n236_));
  XOR2_X1   g035(.A(G71gat), .B(G78gat), .Z(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT12), .B1(new_n233_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(new_n241_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n240_), .B(new_n221_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n245_), .B2(KEYINPUT12), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G230gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT64), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  INV_X1    g051(.A(new_n248_), .ZN(new_n253_));
  NOR4_X1   g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .A4(new_n242_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G120gat), .B(G148gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT5), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n256_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n202_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G15gat), .B(G22gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT75), .B(G8gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G1gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n274_), .B2(KEYINPUT14), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n275_), .A2(new_n276_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(KEYINPUT14), .ZN(new_n283_));
  INV_X1    g082(.A(new_n272_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT76), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n280_), .B1(new_n286_), .B2(new_n277_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G43gat), .B(G50gat), .ZN(new_n289_));
  INV_X1    g088(.A(G36gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G29gat), .ZN(new_n291_));
  INV_X1    g090(.A(G29gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G36gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT71), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n289_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n298_), .A3(new_n289_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(KEYINPUT15), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT15), .ZN(new_n303_));
  INV_X1    g102(.A(new_n301_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n288_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G229gat), .A2(G233gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT79), .Z(new_n309_));
  OAI21_X1  g108(.A(new_n281_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n286_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n304_), .A2(new_n299_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT78), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n315_));
  INV_X1    g114(.A(new_n313_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n315_), .B(new_n316_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n307_), .B(new_n309_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n315_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(KEYINPUT78), .A3(new_n313_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n320_), .A2(new_n321_), .B1(new_n316_), .B2(new_n288_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n318_), .B1(new_n322_), .B2(new_n308_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G113gat), .B(G141gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT80), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G169gat), .B(G197gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n318_), .B(new_n329_), .C1(new_n322_), .C2(new_n308_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n271_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G22gat), .B(G50gat), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G155gat), .B(G162gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G141gat), .B(G148gat), .Z(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n348_), .B(new_n349_), .C1(KEYINPUT1), .C2(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT29), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n352_), .A2(new_n354_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n335_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n357_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n334_), .A3(new_n355_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n360_), .A3(KEYINPUT85), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(G204gat), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G197gat), .A2(G204gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT21), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G218gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G211gat), .ZN(new_n375_));
  INV_X1    g174(.A(G211gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G218gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n367_), .ZN(new_n379_));
  INV_X1    g178(.A(G204gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n372_), .B1(G197gat), .B2(G204gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n373_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n372_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(KEYINPUT88), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT87), .B(G197gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n369_), .B1(new_n390_), .B2(G204gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(new_n386_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n385_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT89), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(KEYINPUT88), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n389_), .A3(new_n386_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n395_), .A2(new_n396_), .B1(new_n373_), .B2(new_n384_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT86), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n351_), .A2(KEYINPUT29), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n394_), .A2(new_n399_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n393_), .A2(new_n402_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n401_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT90), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n403_), .A2(KEYINPUT90), .A3(new_n405_), .A4(new_n408_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n403_), .A2(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n404_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n365_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n365_), .A2(new_n415_), .A3(KEYINPUT91), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(new_n409_), .A3(new_n361_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT25), .B(G183gat), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT81), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G190gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(G183gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT23), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G183gat), .A3(G190gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT23), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT82), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n432_), .B2(KEYINPUT23), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OR3_X1    g240(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n429_), .A2(new_n437_), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G169gat), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n433_), .A2(new_n431_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(G183gat), .A2(G190gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n394_), .A2(new_n399_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT94), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n394_), .A2(new_n399_), .A3(new_n451_), .A4(KEYINPUT94), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G176gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT22), .B(G169gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT93), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n449_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n437_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n464_), .A3(new_n438_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n425_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(new_n423_), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n467_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n397_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(KEYINPUT20), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n456_), .A2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G8gat), .B(G36gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT96), .ZN(new_n478_));
  XOR2_X1   g277(.A(G64gat), .B(G92gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n395_), .A2(new_n396_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n484_), .A2(new_n398_), .A3(new_n385_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n398_), .B1(new_n484_), .B2(new_n385_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n445_), .B(new_n450_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n465_), .A2(new_n468_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n393_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n473_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n476_), .A2(new_n483_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n474_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n482_), .B1(new_n494_), .B2(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT27), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n469_), .A2(KEYINPUT102), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT102), .B1(new_n469_), .B2(new_n498_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n456_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT103), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n472_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n487_), .A2(new_n490_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n473_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n473_), .B1(new_n456_), .B2(new_n501_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n503_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n482_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n493_), .A2(KEYINPUT27), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n496_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G29gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G85gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT0), .B(G57gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G127gat), .B(G134gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G113gat), .B(G120gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n520_), .A2(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n520_), .A2(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(KEYINPUT83), .A3(new_n522_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n351_), .A3(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n347_), .B(new_n350_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(KEYINPUT4), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT97), .B(KEYINPUT4), .Z(new_n534_));
  NAND4_X1  g333(.A1(new_n525_), .A2(new_n351_), .A3(new_n527_), .A4(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n530_), .A2(new_n531_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n528_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n533_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n531_), .B1(new_n540_), .B2(new_n530_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n518_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT104), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n528_), .A2(KEYINPUT4), .A3(new_n529_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT98), .B1(new_n544_), .B2(new_n539_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(new_n517_), .A3(new_n536_), .A4(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT104), .B(new_n518_), .C1(new_n538_), .C2(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G227gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(G15gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT30), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n451_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n525_), .A2(new_n527_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G71gat), .B(G99gat), .ZN(new_n558_));
  INV_X1    g357(.A(G43gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT31), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n557_), .B(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n550_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n422_), .A2(new_n513_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT100), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n538_), .A2(new_n541_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n566_), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n517_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n546_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n528_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n518_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n535_), .A2(new_n532_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n530_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n546_), .B2(new_n569_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n493_), .A2(new_n576_), .A3(new_n495_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n565_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n483_), .B1(new_n476_), .B2(new_n492_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n494_), .A2(new_n482_), .A3(new_n491_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n567_), .A2(new_n570_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n581_), .A2(KEYINPUT100), .A3(new_n582_), .A4(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n509_), .A2(new_n503_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n509_), .A2(new_n503_), .B1(new_n506_), .B2(new_n473_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n492_), .A3(new_n476_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n578_), .B(new_n583_), .C1(new_n587_), .C2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n550_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n590_), .A2(new_n422_), .B1(new_n591_), .B2(new_n513_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n562_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n564_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n333_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n306_), .A2(new_n233_), .A3(KEYINPUT72), .ZN(new_n602_));
  INV_X1    g401(.A(new_n221_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n228_), .A2(new_n230_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT8), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n313_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n599_), .A2(new_n600_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n602_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT72), .B1(new_n306_), .B2(new_n233_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n601_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n607_), .A2(new_n313_), .B1(new_n600_), .B2(new_n599_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n601_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .A4(new_n602_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n596_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT73), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n622_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n617_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  AOI221_X4 g427(.A(new_n596_), .B1(new_n625_), .B2(new_n623_), .C1(new_n612_), .C2(new_n616_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n617_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n612_), .A2(new_n616_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n623_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n634_), .A3(new_n625_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n629_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT37), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n630_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT77), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n312_), .B(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(new_n241_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT16), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n644_), .B(new_n645_), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT17), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n639_), .B1(new_n642_), .B2(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(KEYINPUT17), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n642_), .A2(new_n650_), .A3(new_n648_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n652_), .B1(KEYINPUT77), .B2(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n638_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n595_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(G1gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n550_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(KEYINPUT106), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(KEYINPUT38), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(KEYINPUT106), .A3(new_n659_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n627_), .A2(new_n629_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n653_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n595_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n595_), .A2(KEYINPUT105), .A3(new_n666_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n549_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n662_), .B(new_n663_), .C1(new_n657_), .C2(new_n671_), .ZN(G1324gat));
  INV_X1    g471(.A(new_n513_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n333_), .A2(new_n594_), .A3(new_n673_), .A4(new_n666_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT39), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT107), .B1(new_n674_), .B2(G8gat), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n513_), .A2(new_n273_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n676_), .A2(new_n677_), .B1(new_n656_), .B2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1325gat));
  NAND3_X1  g481(.A1(new_n656_), .A2(new_n552_), .A3(new_n593_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n669_), .A2(new_n670_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n552_), .B1(new_n684_), .B2(new_n593_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT41), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT41), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1326gat));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n422_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n656_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n422_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n689_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n692_), .A2(KEYINPUT42), .A3(new_n689_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(new_n653_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n664_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n595_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n550_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n578_), .A2(new_n583_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n587_), .A2(new_n589_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n422_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n591_), .A2(new_n513_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n593_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n564_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n704_), .B(new_n638_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n704_), .B1(new_n594_), .B2(new_n638_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n333_), .A2(new_n653_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n703_), .B(KEYINPUT44), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n594_), .A2(new_n638_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n703_), .A3(new_n711_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n703_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n549_), .A2(new_n292_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n702_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  NAND4_X1  g524(.A1(new_n595_), .A2(new_n290_), .A3(new_n673_), .A4(new_n699_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n513_), .B1(new_n716_), .B2(new_n722_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n290_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT46), .B(new_n727_), .C1(new_n728_), .C2(new_n290_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  AOI211_X1 g532(.A(new_n559_), .B(new_n562_), .C1(new_n716_), .C2(new_n722_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G43gat), .B1(new_n701_), .B2(new_n593_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT47), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n562_), .A2(new_n559_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n723_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1330gat));
  OR3_X1    g540(.A1(new_n700_), .A2(G50gat), .A3(new_n422_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n723_), .A2(KEYINPUT110), .A3(new_n690_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G50gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT110), .B1(new_n723_), .B2(new_n690_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n742_), .B1(new_n744_), .B2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(G57gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n270_), .A2(new_n331_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n594_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n654_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n750_), .B2(new_n549_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT111), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n666_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n753_), .A2(new_n747_), .A3(new_n549_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n753_), .B2(new_n513_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n513_), .A2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n750_), .B2(new_n759_), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n753_), .B2(new_n562_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n562_), .A2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n750_), .B2(new_n763_), .ZN(G1334gat));
  OR3_X1    g563(.A1(new_n750_), .A2(G78gat), .A3(new_n422_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n749_), .A2(new_n690_), .A3(new_n666_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G78gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT113), .Z(G1335gat));
  NAND2_X1  g570(.A1(new_n749_), .A2(new_n699_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n749_), .A2(new_n774_), .A3(new_n699_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n550_), .ZN(new_n777_));
  NOR4_X1   g576(.A1(new_n714_), .A2(new_n331_), .A3(new_n270_), .A4(new_n698_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n550_), .A2(G85gat), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT115), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(new_n778_), .B2(new_n780_), .ZN(G1336gat));
  NAND3_X1  g580(.A1(new_n776_), .A2(new_n204_), .A3(new_n673_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n778_), .A2(new_n673_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n204_), .ZN(G1337gat));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n209_), .A3(new_n593_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n778_), .A2(new_n593_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n785_), .B(new_n786_), .C1(new_n787_), .C2(new_n223_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n223_), .B1(new_n778_), .B2(new_n593_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n786_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT51), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n791_), .ZN(G1338gat));
  XNOR2_X1  g591(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n270_), .A2(new_n331_), .A3(new_n698_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n690_), .B(new_n795_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(G106gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT52), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n796_), .B2(G106gat), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n776_), .A2(new_n210_), .A3(new_n690_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(G106gat), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(KEYINPUT116), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n794_), .B1(new_n801_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n800_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT52), .A3(new_n798_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(new_n805_), .A3(new_n802_), .A4(new_n793_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1339gat));
  XNOR2_X1  g610(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n628_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n635_), .A2(new_n636_), .A3(KEYINPUT37), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n698_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n269_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n332_), .B1(new_n817_), .B2(new_n265_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n812_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n812_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n654_), .A2(new_n332_), .A3(new_n270_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n331_), .A2(new_n264_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n249_), .A2(new_n254_), .A3(KEYINPUT55), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n246_), .A2(KEYINPUT55), .A3(new_n248_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n253_), .B1(new_n251_), .B2(new_n242_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n261_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n245_), .A2(KEYINPUT12), .ZN(new_n831_));
  INV_X1    g630(.A(new_n242_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n248_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n252_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n246_), .A2(KEYINPUT68), .A3(new_n248_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n825_), .A2(new_n826_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT56), .A3(new_n261_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n823_), .B1(new_n830_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n309_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n307_), .B(new_n842_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n327_), .C1(new_n322_), .C2(new_n842_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n330_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n664_), .B1(new_n841_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n331_), .A2(new_n264_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n839_), .B2(new_n261_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n829_), .B(new_n263_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n262_), .A2(new_n264_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n845_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT57), .A3(new_n664_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n845_), .A2(new_n264_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n830_), .B2(new_n840_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n859_), .B(new_n638_), .C1(new_n861_), .C2(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(KEYINPUT58), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n845_), .A2(new_n264_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n859_), .B1(new_n868_), .B2(new_n638_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n850_), .B(new_n858_), .C1(new_n864_), .C2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n822_), .B1(new_n870_), .B2(new_n653_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n690_), .A2(new_n673_), .A3(new_n549_), .A4(new_n562_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n331_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n815_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n879_), .A2(new_n859_), .B1(KEYINPUT58), .B2(new_n861_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n868_), .A2(new_n638_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT119), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n857_), .B2(new_n664_), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n849_), .B(new_n665_), .C1(new_n854_), .C2(new_n856_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n698_), .B1(new_n883_), .B2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT59), .B(new_n872_), .C1(new_n887_), .C2(new_n822_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n332_), .B1(new_n878_), .B2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n876_), .B1(new_n889_), .B2(new_n875_), .ZN(G1340gat));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n878_), .A2(new_n888_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n271_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n874_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n892_), .B1(new_n270_), .B2(KEYINPUT60), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n892_), .B2(KEYINPUT60), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT120), .B2(new_n896_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n895_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n891_), .B1(new_n894_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n270_), .B1(new_n878_), .B2(new_n888_), .ZN(new_n903_));
  OAI221_X1 g702(.A(KEYINPUT121), .B1(new_n895_), .B2(new_n900_), .C1(new_n903_), .C2(new_n892_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n874_), .A2(new_n906_), .A3(new_n698_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n653_), .B1(new_n878_), .B2(new_n888_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(G1342gat));
  AOI21_X1  g708(.A(G134gat), .B1(new_n874_), .B2(new_n665_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT122), .B(G134gat), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n815_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n893_), .B2(new_n912_), .ZN(G1343gat));
  NOR4_X1   g712(.A1(new_n673_), .A2(new_n422_), .A3(new_n549_), .A4(new_n593_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT123), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n887_), .B2(new_n822_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n332_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT124), .B(G141gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1344gat));
  NOR2_X1   g718(.A1(new_n916_), .A2(new_n270_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n338_), .ZN(G1345gat));
  NOR2_X1   g720(.A1(new_n916_), .A2(new_n653_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT61), .B(G155gat), .Z(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n916_), .B2(new_n815_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n664_), .A2(G162gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n916_), .B2(new_n926_), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n871_), .A2(new_n513_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n422_), .A2(new_n563_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n331_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n932_), .A3(G169gat), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n931_), .B2(G169gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n928_), .A2(new_n930_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n460_), .A2(new_n461_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n332_), .A2(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT125), .ZN(new_n939_));
  OAI22_X1  g738(.A1(new_n934_), .A2(new_n935_), .B1(new_n936_), .B2(new_n939_), .ZN(G1348gat));
  NOR2_X1   g739(.A1(new_n936_), .A2(new_n270_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n457_), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n936_), .A2(new_n653_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(G183gat), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n423_), .B2(new_n943_), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n936_), .B2(new_n815_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n665_), .A2(new_n425_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n936_), .B2(new_n947_), .ZN(G1351gat));
  NAND3_X1  g747(.A1(new_n928_), .A2(new_n591_), .A3(new_n562_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n332_), .ZN(new_n950_));
  INV_X1    g749(.A(G197gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n949_), .A2(new_n270_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT126), .B(G204gat), .Z(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1353gat));
  OAI22_X1  g754(.A1(new_n949_), .A2(new_n653_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n956_));
  OR2_X1    g755(.A1(new_n949_), .A2(new_n653_), .ZN(new_n957_));
  XOR2_X1   g756(.A(KEYINPUT63), .B(G211gat), .Z(new_n958_));
  OAI21_X1  g757(.A(new_n956_), .B1(new_n957_), .B2(new_n958_), .ZN(G1354gat));
  NOR3_X1   g758(.A1(new_n949_), .A2(new_n374_), .A3(new_n815_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n591_), .A2(new_n562_), .ZN(new_n961_));
  NOR4_X1   g760(.A1(new_n871_), .A2(new_n513_), .A3(new_n664_), .A4(new_n961_), .ZN(new_n962_));
  OR2_X1    g761(.A1(new_n962_), .A2(KEYINPUT127), .ZN(new_n963_));
  AOI21_X1  g762(.A(G218gat), .B1(new_n962_), .B2(KEYINPUT127), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n960_), .B1(new_n963_), .B2(new_n964_), .ZN(G1355gat));
endmodule


