//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n211_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n214_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(KEYINPUT84), .A3(new_n212_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219_));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n216_), .B1(new_n213_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n224_), .A2(new_n227_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n225_), .B(new_n226_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n235_), .A2(KEYINPUT90), .A3(new_n218_), .A4(new_n223_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT91), .B1(new_n239_), .B2(KEYINPUT4), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241_));
  AOI211_X1 g040(.A(new_n241_), .B(new_n228_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n232_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n230_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G1gat), .B(G29gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G85gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G57gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  AND3_X1   g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G197gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT86), .B1(new_n254_), .B2(G204gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT86), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(G197gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(G204gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(G197gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT21), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n251_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n255_), .A2(new_n258_), .A3(new_n252_), .A4(new_n259_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n261_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT87), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G218gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G211gat), .ZN(new_n272_));
  INV_X1    g071(.A(G211gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G218gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(KEYINPUT21), .B2(new_n263_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n276_), .A2(new_n266_), .B1(new_n260_), .B2(new_n253_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT87), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n281_), .A2(new_n282_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n287_));
  XOR2_X1   g086(.A(G22gat), .B(G50gat), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n218_), .A2(new_n223_), .A3(new_n290_), .A4(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n287_), .B2(new_n291_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT88), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n287_), .A2(new_n291_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n288_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n300_), .B2(new_n292_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n284_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n300_), .B(new_n292_), .C1(KEYINPUT88), .C2(new_n296_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n281_), .A2(new_n282_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n283_), .A2(new_n280_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n295_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n303_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n249_), .A2(new_n250_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G8gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G169gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(new_n319_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n318_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(KEYINPUT23), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n320_), .A2(KEYINPUT82), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n319_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n319_), .A2(KEYINPUT23), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n326_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G183gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT25), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G183gat), .ZN(new_n337_));
  INV_X1    g136(.A(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT26), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT26), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G190gat), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n335_), .A2(new_n337_), .A3(new_n339_), .A4(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G169gat), .ZN(new_n343_));
  INV_X1    g142(.A(G176gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT24), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(KEYINPUT81), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n333_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT25), .B(G183gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT26), .B(G190gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(G169gat), .B2(G176gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n350_), .A2(new_n351_), .B1(new_n353_), .B2(new_n345_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT81), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n325_), .B1(new_n349_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n316_), .B1(new_n356_), .B2(new_n268_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n324_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n318_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n342_), .A2(new_n347_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n326_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n321_), .C1(new_n322_), .C2(new_n319_), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n361_), .A2(new_n362_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n357_), .B(new_n360_), .C1(new_n268_), .C2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n316_), .B1(new_n366_), .B2(new_n268_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n277_), .B(new_n325_), .C1(new_n349_), .C2(new_n355_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT89), .B1(new_n370_), .B2(new_n359_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n372_));
  AOI211_X1 g171(.A(new_n372_), .B(new_n360_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n315_), .B(new_n367_), .C1(new_n371_), .C2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n320_), .A2(KEYINPUT82), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n327_), .A2(KEYINPUT23), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n319_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n321_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n326_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n324_), .ZN(new_n380_));
  AND2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n382_), .B2(new_n331_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n354_), .A2(new_n379_), .B1(new_n383_), .B2(new_n318_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n270_), .A2(new_n278_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n360_), .B1(new_n357_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n370_), .A2(new_n359_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n374_), .B(KEYINPUT27), .C1(new_n315_), .C2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT92), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n367_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n314_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n374_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI211_X1 g194(.A(KEYINPUT92), .B(KEYINPUT27), .C1(new_n392_), .C2(new_n374_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n310_), .B(new_n389_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n363_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n348_), .A3(new_n333_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n402_), .A2(new_n325_), .A3(new_n277_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n277_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n359_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n372_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n370_), .A2(KEYINPUT89), .A3(new_n359_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n315_), .B1(new_n408_), .B2(new_n367_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n374_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n394_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT92), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n393_), .A2(new_n390_), .A3(new_n394_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n414_), .A2(KEYINPUT93), .A3(new_n310_), .A4(new_n389_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n409_), .A2(new_n410_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n243_), .A2(KEYINPUT33), .A3(new_n244_), .A4(new_n248_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n230_), .B(new_n229_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n248_), .B1(new_n239_), .B2(new_n231_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AND4_X1   g222(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .A4(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n249_), .A2(new_n250_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n315_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(new_n367_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n388_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n309_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n399_), .A2(new_n415_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(G71gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G99gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n356_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(new_n227_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G15gat), .B(G43gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT83), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT30), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT31), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n309_), .B(new_n389_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT94), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n414_), .A2(new_n448_), .A3(new_n309_), .A4(new_n389_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n425_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n445_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n431_), .A2(new_n445_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G29gat), .B(G36gat), .Z(new_n454_));
  XOR2_X1   g253(.A(G43gat), .B(G50gat), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G29gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G43gat), .B(G50gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT15), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G8gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n460_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n460_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n468_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G141gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT80), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G169gat), .B(G197gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n453_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G64gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G57gat), .ZN(new_n490_));
  INV_X1    g289(.A(G57gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G64gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT11), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT69), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G57gat), .B(G64gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT69), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n494_), .ZN(new_n501_));
  AND2_X1   g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT11), .B1(new_n490_), .B2(new_n492_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n506_), .A2(KEYINPUT68), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n499_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT68), .B1(new_n506_), .B2(new_n507_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n504_), .B(new_n500_), .C1(new_n496_), .C2(KEYINPUT11), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n510_), .A2(new_n495_), .A3(new_n498_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(new_n470_), .ZN(new_n514_));
  AND2_X1   g313(.A1(G231gat), .A2(G233gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT16), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n518_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n519_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n519_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n516_), .B(new_n517_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT79), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT79), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n535_));
  AND2_X1   g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G85gat), .ZN(new_n539_));
  INV_X1    g338(.A(G92gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(KEYINPUT67), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT6), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(G99gat), .A3(G106gat), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551_));
  INV_X1    g350(.A(G99gat), .ZN(new_n552_));
  INV_X1    g351(.A(G106gat), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n538_), .A2(new_n543_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n534_), .B(new_n545_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT10), .B(G99gat), .Z(new_n560_));
  AOI22_X1  g359(.A1(new_n560_), .A2(new_n553_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT64), .B(G85gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT65), .B(G92gat), .Z(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT9), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n537_), .B1(new_n536_), .B2(KEYINPUT9), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n561_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n538_), .A2(new_n543_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n547_), .A2(new_n549_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n555_), .A3(new_n554_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n569_), .B(new_n571_), .C1(new_n544_), .C2(KEYINPUT8), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n559_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT75), .B1(new_n461_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n573_), .A2(KEYINPUT74), .A3(new_n474_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT74), .B1(new_n573_), .B2(new_n474_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n461_), .A2(new_n573_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G190gat), .B(G218gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT76), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n580_), .A2(new_n582_), .A3(new_n581_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n574_), .A2(new_n578_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT77), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n585_), .A2(KEYINPUT77), .A3(new_n591_), .A4(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n589_), .B(new_n590_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n585_), .B2(new_n594_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n533_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n533_), .ZN(new_n604_));
  AOI211_X1 g403(.A(new_n601_), .B(new_n604_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n532_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n545_), .A2(new_n534_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n569_), .A2(new_n571_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT65), .B(G92gat), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n562_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n566_), .B1(new_n611_), .B2(KEYINPUT9), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n608_), .A2(new_n609_), .B1(new_n612_), .B2(new_n561_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n613_), .A2(new_n512_), .A3(new_n509_), .A4(new_n572_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n573_), .A2(new_n513_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n607_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT70), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n573_), .A2(new_n513_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n607_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT70), .B(new_n607_), .C1(new_n573_), .C2(new_n513_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n573_), .A2(new_n513_), .A3(KEYINPUT12), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT12), .B1(new_n573_), .B2(new_n513_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n616_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT5), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT71), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n626_), .A2(KEYINPUT72), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT72), .B1(new_n626_), .B2(new_n632_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n630_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT13), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n633_), .B(new_n639_), .C1(new_n636_), .C2(new_n634_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n606_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n488_), .A2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(G1gat), .A3(new_n425_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT38), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT38), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n601_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n453_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n532_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n641_), .A2(new_n487_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n425_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n646_), .A3(new_n652_), .ZN(G1324gat));
  NAND2_X1  g452(.A1(new_n414_), .A2(new_n389_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n464_), .A2(new_n488_), .A3(new_n654_), .A4(new_n642_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT95), .ZN(new_n656_));
  INV_X1    g455(.A(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n651_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n656_), .A2(new_n660_), .A3(KEYINPUT40), .A4(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  OAI21_X1  g465(.A(G15gat), .B1(new_n651_), .B2(new_n445_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT41), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n643_), .A2(G15gat), .A3(new_n445_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1326gat));
  XNOR2_X1  g469(.A(new_n309_), .B(KEYINPUT96), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n643_), .A2(G22gat), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n648_), .A2(new_n650_), .A3(new_n671_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(G22gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n674_), .B2(G22gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n673_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT97), .Z(G1327gat));
  INV_X1    g479(.A(new_n641_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n647_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n532_), .A2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT99), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n488_), .A2(new_n681_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n451_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n641_), .A2(new_n487_), .A3(new_n532_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n431_), .A2(new_n445_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n450_), .A2(new_n452_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n647_), .B(new_n533_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n689_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT43), .B(new_n693_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n688_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(KEYINPUT98), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT98), .ZN(new_n700_));
  INV_X1    g499(.A(new_n688_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n453_), .B2(new_n693_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .A4(new_n423_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n309_), .A2(new_n704_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n444_), .B1(new_n705_), .B2(new_n415_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n452_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n689_), .B(new_n694_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n701_), .B1(new_n702_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n700_), .B1(new_n710_), .B2(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n699_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT44), .B(new_n688_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n451_), .A2(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n687_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n654_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n712_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n654_), .A2(new_n719_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n685_), .A2(KEYINPUT45), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT45), .B1(new_n685_), .B2(new_n723_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n718_), .B1(new_n722_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n720_), .B1(new_n711_), .B2(new_n699_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT46), .B(new_n726_), .C1(new_n729_), .C2(new_n719_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1329gat));
  AOI211_X1 g530(.A(new_n698_), .B(new_n701_), .C1(new_n702_), .C2(new_n709_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n444_), .A2(G43gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n732_), .B(new_n733_), .C1(new_n699_), .C2(new_n711_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G43gat), .B1(new_n686_), .B2(new_n444_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT47), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(new_n735_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n737_), .B(new_n738_), .C1(new_n714_), .C2(new_n733_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n686_), .B2(new_n671_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n309_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n715_), .B2(new_n743_), .ZN(G1331gat));
  NAND4_X1  g543(.A1(new_n648_), .A2(new_n487_), .A3(new_n641_), .A4(new_n532_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n425_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n641_), .A2(new_n487_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n453_), .A2(new_n606_), .A3(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n491_), .A3(new_n451_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT100), .ZN(G1332gat));
  OAI21_X1  g550(.A(G64gat), .B1(new_n745_), .B2(new_n657_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT48), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n489_), .A3(new_n654_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n433_), .A3(new_n444_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G71gat), .B1(new_n745_), .B2(new_n445_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT102), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT102), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT101), .B(KEYINPUT49), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n761_), .B2(new_n762_), .ZN(G1334gat));
  OAI21_X1  g562(.A(G78gat), .B1(new_n745_), .B2(new_n672_), .ZN(new_n764_));
  XOR2_X1   g563(.A(KEYINPUT103), .B(KEYINPUT50), .Z(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(G78gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n748_), .A2(new_n767_), .A3(new_n671_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1335gat));
  NAND3_X1  g568(.A1(new_n641_), .A2(new_n487_), .A3(new_n649_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT104), .Z(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n702_), .B2(new_n709_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n451_), .A3(new_n563_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n453_), .A2(new_n747_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n684_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n539_), .B1(new_n775_), .B2(new_n425_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT105), .ZN(G1336gat));
  OAI21_X1  g577(.A(new_n540_), .B1(new_n775_), .B2(new_n657_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT106), .Z(new_n780_));
  NAND2_X1  g579(.A1(new_n654_), .A2(new_n564_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT107), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n772_), .B2(new_n782_), .ZN(G1337gat));
  AOI21_X1  g582(.A(new_n552_), .B1(new_n772_), .B2(new_n444_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n775_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n444_), .A2(new_n560_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n553_), .A3(new_n742_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n772_), .A2(new_n742_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G106gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT52), .B(new_n553_), .C1(new_n772_), .C2(new_n742_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n790_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n642_), .B2(new_n487_), .ZN(new_n801_));
  NOR4_X1   g600(.A1(new_n606_), .A2(new_n641_), .A3(KEYINPUT54), .A4(new_n486_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n469_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n475_), .A2(new_n472_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n483_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n485_), .B1(new_n806_), .B2(KEYINPUT111), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(KEYINPUT111), .B2(new_n806_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n633_), .B(new_n808_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n635_), .A2(new_n486_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT70), .B1(new_n614_), .B2(new_n607_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n621_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n625_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n622_), .A2(KEYINPUT55), .A3(new_n625_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n625_), .A2(new_n614_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n619_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n631_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT109), .B(KEYINPUT56), .Z(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n631_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n810_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n809_), .B1(new_n825_), .B2(KEYINPUT110), .ZN(new_n826_));
  INV_X1    g625(.A(new_n810_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n824_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n821_), .B1(new_n819_), .B2(new_n631_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(KEYINPUT110), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n682_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n808_), .A2(new_n635_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT112), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n808_), .A2(new_n837_), .A3(new_n635_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n631_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n824_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT113), .B(KEYINPUT56), .C1(new_n819_), .C2(new_n631_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n693_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n839_), .B(KEYINPUT58), .C1(new_n842_), .C2(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT57), .B(new_n682_), .C1(new_n826_), .C2(new_n831_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n834_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n803_), .B1(new_n850_), .B2(new_n649_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n450_), .A2(new_n444_), .A3(new_n451_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n851_), .A2(new_n487_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G113gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(KEYINPUT114), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n853_), .B2(G113gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n852_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861_));
  INV_X1    g660(.A(new_n852_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n863_));
  AOI22_X1  g662(.A1(new_n832_), .A2(new_n833_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n532_), .B1(new_n864_), .B2(new_n849_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n862_), .B(new_n863_), .C1(new_n865_), .C2(new_n803_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n860_), .A2(new_n861_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n861_), .B1(new_n860_), .B2(new_n866_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n487_), .A2(new_n855_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n859_), .B1(new_n869_), .B2(new_n870_), .ZN(G1340gat));
  NOR2_X1   g670(.A1(new_n851_), .A2(new_n852_), .ZN(new_n872_));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n681_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n872_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n873_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n860_), .A2(new_n866_), .A3(new_n641_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT117), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G120gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(KEYINPUT117), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n872_), .B2(new_n532_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n649_), .A2(KEYINPUT118), .ZN(new_n882_));
  MUX2_X1   g681(.A(KEYINPUT118), .B(new_n882_), .S(G127gat), .Z(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n869_), .B2(new_n883_), .ZN(G1342gat));
  INV_X1    g683(.A(G134gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n872_), .A2(new_n885_), .A3(new_n647_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n867_), .A2(new_n868_), .A3(new_n693_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1343gat));
  NAND4_X1  g687(.A1(new_n657_), .A2(new_n445_), .A3(new_n451_), .A4(new_n742_), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n851_), .A2(KEYINPUT119), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n851_), .B2(new_n889_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n487_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT120), .B(G141gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1344gat));
  AOI21_X1  g693(.A(new_n681_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT121), .B(G148gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1345gat));
  AOI21_X1  g696(.A(new_n649_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n898_), .B(new_n900_), .ZN(G1346gat));
  NAND2_X1  g700(.A1(new_n890_), .A2(new_n891_), .ZN(new_n902_));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n647_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n693_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1347gat));
  NOR2_X1   g705(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n657_), .A2(new_n707_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n672_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n851_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(KEYINPUT123), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n851_), .A2(new_n913_), .A3(new_n910_), .ZN(new_n914_));
  OAI221_X1 g713(.A(new_n486_), .B1(new_n907_), .B2(new_n908_), .C1(new_n912_), .C2(new_n914_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n851_), .A2(new_n487_), .A3(new_n910_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n343_), .B1(new_n916_), .B2(KEYINPUT122), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  INV_X1    g717(.A(new_n910_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n486_), .B(new_n919_), .C1(new_n865_), .C2(new_n803_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n917_), .A2(new_n918_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n918_), .B1(new_n917_), .B2(new_n922_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n915_), .B1(new_n923_), .B2(new_n924_), .ZN(G1348gat));
  OAI21_X1  g724(.A(new_n641_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n851_), .A2(new_n742_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n681_), .A2(new_n657_), .A3(new_n344_), .A4(new_n707_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n926_), .A2(new_n344_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  INV_X1    g728(.A(new_n912_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n914_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n649_), .A2(new_n350_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n927_), .A2(new_n532_), .A3(new_n909_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n932_), .A2(new_n933_), .B1(new_n334_), .B2(new_n934_), .ZN(G1350gat));
  OAI211_X1 g734(.A(new_n351_), .B(new_n647_), .C1(new_n912_), .C2(new_n914_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n693_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n338_), .ZN(G1351gat));
  NAND3_X1  g737(.A1(new_n654_), .A2(new_n445_), .A3(new_n310_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n851_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n486_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g741(.A1(new_n851_), .A2(new_n681_), .A3(new_n939_), .ZN(new_n943_));
  AND2_X1   g742(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n945_), .ZN(G1353gat));
  AOI21_X1  g746(.A(new_n649_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n948_));
  XOR2_X1   g747(.A(new_n948_), .B(KEYINPUT125), .Z(new_n949_));
  NAND2_X1  g748(.A1(new_n940_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  XOR2_X1   g750(.A(new_n950_), .B(new_n951_), .Z(G1354gat));
  AOI21_X1  g751(.A(G218gat), .B1(new_n940_), .B2(new_n647_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n693_), .A2(new_n271_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT126), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n940_), .B2(new_n955_), .ZN(G1355gat));
endmodule


