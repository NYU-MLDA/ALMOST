//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  XOR2_X1   g000(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n212_), .B(new_n213_), .C1(new_n214_), .C2(new_n210_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n221_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n215_), .A2(new_n220_), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n223_), .A3(KEYINPUT83), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n224_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n229_));
  OR2_X1    g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n219_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(new_n217_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT21), .B1(new_n236_), .B2(KEYINPUT87), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  INV_X1    g037(.A(G218gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(G211gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(G211gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G197gat), .B(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n237_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(KEYINPUT21), .B(new_n243_), .C1(new_n236_), .C2(KEYINPUT87), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n227_), .A2(new_n235_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n247_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT90), .B1(new_n247_), .B2(KEYINPUT20), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n246_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n225_), .A2(new_n223_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n230_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n234_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n214_), .A2(new_n213_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n220_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n221_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n228_), .A2(new_n229_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT91), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n228_), .A2(new_n229_), .A3(new_n260_), .A4(new_n257_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n256_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n254_), .B1(new_n262_), .B2(KEYINPUT92), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT92), .ZN(new_n264_));
  AOI211_X1 g063(.A(new_n264_), .B(new_n256_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n251_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n209_), .B1(new_n250_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n227_), .A2(new_n235_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n251_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(KEYINPUT20), .A3(new_n209_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n263_), .A2(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n251_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n206_), .B1(new_n267_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT94), .B(new_n206_), .C1(new_n267_), .C2(new_n273_), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n267_), .A2(new_n273_), .A3(new_n206_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n250_), .A2(new_n209_), .A3(new_n266_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n272_), .A2(new_n254_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(new_n262_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n269_), .A2(KEYINPUT20), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n208_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n206_), .B(KEYINPUT97), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n278_), .A2(KEYINPUT27), .A3(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n281_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G113gat), .B(G120gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G155gat), .B(G162gat), .ZN(new_n298_));
  INV_X1    g097(.A(G141gat), .ZN(new_n299_));
  INV_X1    g098(.A(G148gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT3), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(G141gat), .B2(G148gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n298_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G155gat), .B(G162gat), .Z(new_n313_));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n296_), .B(new_n297_), .C1(new_n308_), .C2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n292_), .A2(new_n293_), .ZN(new_n319_));
  INV_X1    g118(.A(G127gat), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n320_), .A2(G134gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(G134gat), .ZN(new_n322_));
  INV_X1    g121(.A(G113gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(G120gat), .ZN(new_n324_));
  INV_X1    g123(.A(G120gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(G113gat), .ZN(new_n326_));
  OAI22_X1  g125(.A1(new_n321_), .A2(new_n322_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n319_), .B(new_n327_), .C1(new_n315_), .C2(new_n308_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n304_), .A2(new_n307_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n313_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n309_), .A2(new_n310_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n331_), .B(new_n311_), .C1(KEYINPUT1), .C2(new_n298_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n319_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n334_), .A3(KEYINPUT4), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n332_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(KEYINPUT95), .A3(new_n297_), .A4(new_n296_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n318_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT0), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G57gat), .ZN(new_n348_));
  INV_X1    g147(.A(G85gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n342_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n268_), .B(KEYINPUT30), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT84), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n357_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(new_n296_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT31), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n362_), .B(new_n333_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n365_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n251_), .B2(KEYINPUT88), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n336_), .A2(KEYINPUT29), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT89), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n251_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n379_), .B2(new_n251_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n378_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n378_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n336_), .A2(KEYINPUT29), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT28), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n385_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n291_), .A2(new_n356_), .A3(new_n371_), .A4(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT100), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT99), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n318_), .A2(new_n335_), .A3(new_n339_), .A4(new_n337_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n328_), .A2(new_n340_), .A3(new_n334_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n350_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n344_), .A2(new_n405_), .A3(new_n351_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT33), .B1(new_n353_), .B2(new_n350_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n276_), .A2(new_n408_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT32), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n206_), .A2(new_n410_), .ZN(new_n411_));
  OR3_X1    g210(.A1(new_n267_), .A2(new_n273_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n287_), .A2(new_n411_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n355_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n398_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT96), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT98), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n279_), .A2(new_n280_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n398_), .A2(new_n355_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n290_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT96), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n415_), .A2(new_n423_), .A3(new_n398_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n281_), .A2(KEYINPUT98), .A3(new_n420_), .A4(new_n290_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n417_), .A2(new_n422_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n370_), .B(KEYINPUT85), .Z(new_n427_));
  AOI21_X1  g226(.A(new_n401_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n401_), .A3(new_n427_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n400_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT12), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G57gat), .B(G64gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT11), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G78gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n438_), .B(new_n439_), .C1(KEYINPUT11), .C2(new_n433_), .ZN(new_n440_));
  INV_X1    g239(.A(G64gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G57gat), .ZN(new_n442_));
  INV_X1    g241(.A(G57gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G64gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT11), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT67), .B1(new_n445_), .B2(new_n437_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n440_), .A2(new_n446_), .A3(new_n436_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(KEYINPUT71), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT71), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n440_), .A2(new_n446_), .A3(new_n436_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n447_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n432_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT65), .B(G85gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n460_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT64), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT64), .ZN(new_n474_));
  NOR4_X1   g273(.A1(new_n469_), .A2(new_n470_), .A3(new_n474_), .A4(G106gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n455_), .B1(new_n468_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT10), .B(G99gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n474_), .B1(new_n478_), .B2(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(KEYINPUT64), .A3(new_n472_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G92gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI22_X1  g284(.A1(new_n485_), .A2(new_n462_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n481_), .A2(new_n486_), .A3(KEYINPUT69), .A4(new_n460_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n477_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n489_));
  INV_X1    g288(.A(G99gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n472_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n491_), .A2(new_n458_), .A3(new_n459_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n349_), .A2(new_n482_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n465_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT68), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT8), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n488_), .A2(new_n506_), .A3(KEYINPUT70), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT70), .B1(new_n488_), .B2(new_n506_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n454_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n452_), .A2(new_n447_), .ZN(new_n511_));
  OAI22_X1  g310(.A1(new_n468_), .A2(new_n476_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT12), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n511_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n514_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(G230gat), .A3(G233gat), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G176gat), .B(G204gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G120gat), .B(G148gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT73), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n525_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n528_), .B(KEYINPUT74), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n522_), .A2(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n530_), .A2(new_n533_), .A3(KEYINPUT13), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT13), .B1(new_n530_), .B2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT77), .B(G15gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(G22gat), .ZN(new_n538_));
  INV_X1    g337(.A(G1gat), .ZN(new_n539_));
  INV_X1    g338(.A(G8gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT14), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT78), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n544_), .A3(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G1gat), .B(G8gat), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n547_), .A3(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G43gat), .B(G50gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT76), .ZN(new_n554_));
  INV_X1    g353(.A(G29gat), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G36gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(G36gat), .A3(new_n557_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n560_), .A2(KEYINPUT15), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT15), .B1(new_n560_), .B2(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n552_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n561_), .ZN(new_n566_));
  AOI21_X1  g365(.A(G36gat), .B1(new_n556_), .B2(new_n557_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT81), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n551_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n551_), .B2(new_n568_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n564_), .B(new_n565_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n551_), .A2(new_n568_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n551_), .A2(new_n568_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT81), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n576_), .B2(new_n570_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n573_), .B1(new_n577_), .B2(new_n565_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(G169gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(G197gat), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n573_), .B(new_n581_), .C1(new_n577_), .C2(new_n565_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n536_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT34), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n590_));
  AOI22_X1  g389(.A1(new_n568_), .A2(new_n518_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n562_), .A2(new_n563_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n507_), .A2(new_n508_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(new_n590_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n595_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n596_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n599_), .B(KEYINPUT36), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT37), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(KEYINPUT37), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n551_), .B(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n613_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n612_), .A2(new_n511_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n612_), .A2(new_n511_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n619_), .B(new_n614_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT80), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n610_), .A2(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n431_), .A2(new_n586_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n539_), .A3(new_n355_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT38), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n399_), .B(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n426_), .A2(new_n401_), .A3(new_n427_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(new_n428_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n586_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n628_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n606_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n636_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n641_), .B2(new_n356_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n632_), .A2(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(new_n291_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n540_), .B1(new_n640_), .B2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT39), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n291_), .A2(G8gat), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n646_), .A2(new_n650_), .B1(new_n630_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1325gat));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n427_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n640_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT102), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n630_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n397_), .B(KEYINPUT103), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n640_), .B2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT42), .Z(new_n667_));
  NAND3_X1  g466(.A1(new_n630_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n606_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n586_), .A2(new_n628_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n431_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n355_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n636_), .A2(new_n675_), .A3(new_n609_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n636_), .B2(new_n609_), .ZN(new_n677_));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n671_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(G29gat), .A3(new_n355_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n676_), .A2(new_n677_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n672_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n674_), .B1(new_n679_), .B2(new_n682_), .ZN(G1328gat));
  AND2_X1   g482(.A1(new_n678_), .A2(new_n644_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n559_), .B1(new_n684_), .B2(new_n682_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n673_), .A2(new_n559_), .A3(new_n644_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT46), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n685_), .A2(new_n688_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n685_), .B2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  NAND3_X1  g492(.A1(new_n678_), .A2(G43gat), .A3(new_n371_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n431_), .B2(new_n610_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n636_), .A2(new_n675_), .A3(new_n609_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n671_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n673_), .A2(new_n657_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT106), .B(G43gat), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n694_), .A2(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g501(.A(G50gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n673_), .A2(new_n703_), .A3(new_n665_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n682_), .A2(new_n397_), .A3(new_n678_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n682_), .A2(KEYINPUT107), .A3(new_n397_), .A4(new_n678_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n678_), .A2(new_n397_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n711_), .B2(new_n698_), .ZN(new_n712_));
  AND4_X1   g511(.A1(new_n705_), .A2(new_n712_), .A3(new_n709_), .A4(G50gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n704_), .B1(new_n710_), .B2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n629_), .A2(new_n536_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT109), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n716_), .A2(new_n585_), .A3(new_n431_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n443_), .A3(new_n355_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n636_), .A2(new_n639_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n536_), .A2(new_n585_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n356_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(G1332gat));
  AOI21_X1  g523(.A(new_n441_), .B1(new_n721_), .B2(new_n644_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT48), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n717_), .A2(new_n441_), .A3(new_n644_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1333gat));
  NOR2_X1   g527(.A1(new_n427_), .A2(G71gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n717_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n721_), .A2(new_n657_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G71gat), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(KEYINPUT110), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(KEYINPUT110), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(KEYINPUT49), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT49), .B1(new_n734_), .B2(new_n735_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n731_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n721_), .B2(new_n665_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT50), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n717_), .A2(new_n739_), .A3(new_n665_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n720_), .A2(new_n638_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n636_), .A2(new_n606_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n355_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n681_), .A2(new_n744_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n355_), .A2(new_n463_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT112), .Z(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n749_), .B2(new_n751_), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n747_), .A2(new_n482_), .A3(new_n644_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n681_), .A2(new_n291_), .A3(new_n744_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n482_), .ZN(G1337gat));
  NAND3_X1  g554(.A1(new_n747_), .A2(new_n471_), .A3(new_n371_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n681_), .A2(new_n427_), .A3(new_n744_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n490_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n747_), .A2(new_n472_), .A3(new_n397_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n397_), .B(new_n745_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n697_), .A2(KEYINPUT113), .A3(new_n397_), .A4(new_n745_), .ZN(new_n765_));
  AND4_X1   g564(.A1(new_n761_), .A2(new_n764_), .A3(G106gat), .A4(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n472_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n761_), .B1(new_n767_), .B2(new_n765_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n760_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n760_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n510_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n516_), .A2(KEYINPUT114), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(KEYINPUT55), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n516_), .A2(KEYINPUT114), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n532_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT56), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n780_), .B2(KEYINPUT56), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n777_), .A2(new_n779_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n531_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n565_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n564_), .B(new_n790_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n582_), .C1(new_n577_), .C2(new_n790_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n584_), .A2(new_n792_), .A3(new_n529_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n774_), .B1(new_n784_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n786_), .A2(new_n788_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT117), .A3(new_n781_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(KEYINPUT58), .A3(new_n789_), .A4(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n609_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n788_), .B1(new_n780_), .B2(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n516_), .A2(KEYINPUT114), .A3(new_n778_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n778_), .B1(new_n516_), .B2(KEYINPUT114), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n775_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT115), .B(KEYINPUT56), .C1(new_n805_), .C2(new_n532_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n530_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n802_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n584_), .B(new_n792_), .C1(new_n530_), .C2(new_n533_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n606_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n800_), .B1(new_n810_), .B2(KEYINPUT116), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n812_), .B(new_n606_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n799_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n638_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n536_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n585_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n610_), .A2(new_n628_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n610_), .A2(new_n819_), .A3(new_n822_), .A4(new_n628_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n817_), .A2(new_n824_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n644_), .A2(new_n356_), .A3(new_n370_), .A4(new_n397_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  INV_X1    g628(.A(new_n824_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n799_), .B(new_n832_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n815_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n830_), .B1(new_n834_), .B2(new_n638_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n826_), .A2(new_n829_), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n828_), .A2(new_n829_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n585_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G113gat), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n828_), .A2(new_n323_), .A3(new_n585_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n837_), .B2(new_n536_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n325_), .A2(KEYINPUT60), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n325_), .B1(new_n536_), .B2(KEYINPUT60), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n845_), .B2(new_n844_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n842_), .B1(new_n827_), .B2(new_n847_), .ZN(G1341gat));
  NAND2_X1  g647(.A1(new_n628_), .A2(G127gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT120), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n837_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n320_), .B1(new_n827_), .B2(new_n638_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n837_), .B2(new_n610_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n670_), .A2(G134gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n827_), .B2(new_n855_), .ZN(G1343gat));
  NOR4_X1   g655(.A1(new_n657_), .A2(new_n356_), .A3(new_n398_), .A4(new_n644_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n825_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n838_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT121), .B(G141gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n858_), .A2(new_n536_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n300_), .ZN(G1345gat));
  NAND3_X1  g662(.A1(new_n825_), .A2(new_n628_), .A3(new_n857_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT122), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n825_), .A2(new_n866_), .A3(new_n628_), .A4(new_n857_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT61), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n870_), .A3(new_n867_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n869_), .A2(G155gat), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G155gat), .B1(new_n869_), .B2(new_n871_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1346gat));
  NOR2_X1   g673(.A1(new_n858_), .A2(new_n670_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n609_), .A2(G162gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT123), .Z(new_n877_));
  OAI22_X1  g676(.A1(new_n875_), .A2(G162gat), .B1(new_n858_), .B2(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT124), .Z(G1347gat));
  NOR3_X1   g678(.A1(new_n427_), .A2(new_n355_), .A3(new_n291_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n665_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n816_), .B1(new_n814_), .B2(KEYINPUT118), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n628_), .B1(new_n883_), .B2(new_n833_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n585_), .B(new_n882_), .C1(new_n884_), .C2(new_n830_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n216_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n882_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT126), .B1(new_n835_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n882_), .C1(new_n884_), .C2(new_n830_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n585_), .A2(new_n233_), .ZN(new_n897_));
  OAI22_X1  g696(.A1(new_n890_), .A2(new_n891_), .B1(new_n896_), .B2(new_n897_), .ZN(G1348gat));
  NAND2_X1  g697(.A1(new_n825_), .A2(new_n398_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n899_), .A2(new_n217_), .A3(new_n536_), .A4(new_n881_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n893_), .A2(new_n818_), .A3(new_n895_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n217_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT127), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n901_), .A2(KEYINPUT127), .A3(new_n217_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n900_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NOR3_X1   g705(.A1(new_n896_), .A2(new_n213_), .A3(new_n638_), .ZN(new_n907_));
  INV_X1    g706(.A(G183gat), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n825_), .A2(new_n398_), .A3(new_n628_), .A4(new_n880_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n896_), .B2(new_n610_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n606_), .A2(new_n214_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n896_), .B2(new_n912_), .ZN(G1351gat));
  AND4_X1   g712(.A1(new_n427_), .A2(new_n825_), .A3(new_n420_), .A4(new_n644_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n585_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n818_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n628_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  NAND3_X1  g722(.A1(new_n914_), .A2(new_n239_), .A3(new_n606_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n914_), .A2(new_n609_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n239_), .ZN(G1355gat));
endmodule


