//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT74), .ZN(new_n203_));
  XOR2_X1   g002(.A(G43gat), .B(G50gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n205_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n205_), .B(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n212_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n205_), .A2(new_n213_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G169gat), .B(G197gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(new_n223_), .A3(new_n227_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n224_), .A2(KEYINPUT81), .A3(new_n228_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(KEYINPUT24), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT23), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT83), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n238_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT25), .B(G183gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT26), .B(G190gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n237_), .A2(KEYINPUT24), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT82), .ZN(new_n252_));
  INV_X1    g051(.A(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT22), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT84), .B1(new_n254_), .B2(G169gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(new_n255_), .C1(new_n256_), .C2(KEYINPUT84), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n240_), .A2(new_n244_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n258_), .A2(new_n260_), .B1(G169gat), .B2(G176gat), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n245_), .A2(new_n252_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(G197gat), .B(G204gat), .Z(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(KEYINPUT21), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n263_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(KEYINPUT21), .ZN(new_n267_));
  MUX2_X1   g066(.A(new_n263_), .B(new_n266_), .S(new_n267_), .Z(new_n268_));
  NOR2_X1   g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n256_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n249_), .B1(new_n275_), .B2(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n242_), .A2(new_n244_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n276_), .B1(new_n277_), .B2(new_n260_), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n236_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n258_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT90), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT90), .B1(new_n280_), .B2(new_n258_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n248_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT89), .ZN(new_n286_));
  INV_X1    g085(.A(new_n249_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n279_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n279_), .B2(new_n287_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n237_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT91), .B1(new_n285_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n281_), .B(new_n282_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n248_), .A4(new_n290_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n278_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n268_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n274_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n270_), .B1(new_n262_), .B2(new_n268_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n296_), .B2(new_n268_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(KEYINPUT92), .A3(new_n273_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT92), .B1(new_n300_), .B2(new_n273_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n298_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G8gat), .B(G36gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT94), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n298_), .B(new_n309_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n304_), .A2(KEYINPUT94), .A3(new_n310_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n278_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n268_), .B(new_n318_), .C1(new_n291_), .C2(new_n285_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n319_), .B(KEYINPUT20), .C1(new_n262_), .C2(new_n268_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n273_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n300_), .B2(new_n273_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n315_), .B1(new_n322_), .B2(new_n310_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n313_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G155gat), .B(G162gat), .Z(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G148gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n328_), .A2(new_n329_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(KEYINPUT85), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n337_), .C1(new_n338_), .C2(KEYINPUT2), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(KEYINPUT2), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n326_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT28), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n342_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n268_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(G78gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G106gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n351_), .B(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n349_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n347_), .A2(new_n348_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n349_), .A2(new_n359_), .A3(new_n357_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n325_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT96), .B(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n342_), .A2(KEYINPUT95), .ZN(new_n369_));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(G113gat), .B(G120gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n369_), .B(new_n372_), .Z(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(KEYINPUT97), .A3(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(KEYINPUT4), .ZN(new_n380_));
  INV_X1    g179(.A(new_n374_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n350_), .A2(new_n382_), .A3(new_n372_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n368_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n368_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(new_n377_), .A3(new_n387_), .A4(new_n378_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(KEYINPUT99), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT99), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n368_), .C1(new_n379_), .C2(new_n384_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G71gat), .B(G99gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G43gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n262_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(new_n372_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(G15gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT30), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT31), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n397_), .A2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n393_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n363_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n379_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n409_), .A2(KEYINPUT33), .A3(new_n387_), .A4(new_n386_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n387_), .B1(new_n373_), .B2(new_n381_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT98), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n380_), .A2(new_n374_), .A3(new_n383_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n412_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n388_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n300_), .A2(new_n273_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT92), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n423_), .A2(new_n301_), .B1(new_n297_), .B2(new_n274_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT32), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n310_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n322_), .A2(KEYINPUT32), .A3(new_n309_), .ZN(new_n427_));
  AND4_X1   g226(.A1(new_n426_), .A2(new_n389_), .A3(new_n391_), .A4(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n361_), .B1(new_n420_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n361_), .B1(new_n391_), .B2(new_n389_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n405_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT100), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n408_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n433_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n235_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G127gat), .B(G155gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT16), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G183gat), .B(G211gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT78), .Z(new_n442_));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n442_), .A2(new_n443_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G231gat), .A2(G233gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n212_), .B(new_n446_), .Z(new_n447_));
  XNOR2_X1  g246(.A(G57gat), .B(G64gat), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n448_), .A2(KEYINPUT11), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(KEYINPUT11), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G71gat), .B(G78gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n448_), .A2(new_n451_), .A3(KEYINPUT11), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n447_), .B(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n444_), .A2(new_n445_), .A3(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT79), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n450_), .A2(new_n452_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n448_), .A2(KEYINPUT11), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n459_), .B(new_n454_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n447_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n447_), .A2(new_n466_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n469_));
  NOR4_X1   g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n441_), .A4(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n458_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT9), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT64), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT10), .B(G99gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(G106gat), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n490_));
  INV_X1    g289(.A(G99gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n355_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT65), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n355_), .A4(KEYINPUT65), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n494_), .A2(new_n486_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n473_), .A2(KEYINPUT66), .A3(new_n475_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT8), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT68), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n489_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n220_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n489_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT67), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT67), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n489_), .B(new_n512_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n205_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT73), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n509_), .A2(new_n515_), .A3(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n521_), .A2(new_n522_), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G190gat), .B(G218gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(G134gat), .B(G162gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n532_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n528_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n526_), .B(new_n527_), .C1(new_n537_), .C2(new_n533_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(KEYINPUT37), .A3(new_n538_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n472_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n455_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n511_), .A2(new_n513_), .A3(new_n544_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT12), .B1(new_n463_), .B2(new_n464_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n508_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n489_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n502_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n505_), .A2(KEYINPUT68), .A3(new_n506_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT70), .B1(new_n556_), .B2(new_n550_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n548_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n545_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n547_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n565_), .A2(new_n571_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(KEYINPUT72), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT72), .B1(new_n573_), .B2(new_n574_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(KEYINPUT13), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n437_), .A2(new_n543_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n207_), .A3(new_n393_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n539_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n580_), .A2(new_n235_), .A3(new_n472_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n589_), .B2(new_n392_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n584_), .A2(new_n585_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n586_), .B(new_n590_), .C1(new_n593_), .C2(new_n594_), .ZN(G1324gat));
  INV_X1    g394(.A(new_n325_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n582_), .A2(G8gat), .A3(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G8gat), .B1(new_n589_), .B2(new_n596_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT39), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT39), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n597_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n601_), .B(new_n603_), .ZN(G1325gat));
  OAI21_X1  g403(.A(G15gat), .B1(new_n589_), .B2(new_n406_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT41), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n583_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  OAI21_X1  g407(.A(G22gat), .B1(new_n589_), .B2(new_n361_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT42), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n361_), .A2(G22gat), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n610_), .B1(new_n582_), .B2(new_n611_), .ZN(G1327gat));
  NOR3_X1   g411(.A1(new_n580_), .A2(new_n235_), .A3(new_n471_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n429_), .A2(new_n431_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n406_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT100), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n436_), .A3(new_n408_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n541_), .A2(new_n542_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n614_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT100), .B(new_n405_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n614_), .B(new_n620_), .C1(new_n434_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n613_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT44), .B(new_n613_), .C1(new_n621_), .C2(new_n624_), .ZN(new_n628_));
  AND4_X1   g427(.A1(G29gat), .A2(new_n627_), .A3(new_n393_), .A4(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630_));
  INV_X1    g429(.A(new_n539_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n580_), .A2(new_n631_), .A3(new_n471_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n234_), .B(new_n632_), .C1(new_n434_), .C2(new_n622_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n393_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n629_), .A2(new_n630_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n630_), .B1(new_n629_), .B2(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1328gat));
  NAND3_X1  g437(.A1(new_n627_), .A2(new_n325_), .A3(new_n628_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G36gat), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n596_), .A2(G36gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT104), .B1(new_n633_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT45), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n647_), .A2(new_n649_), .B1(KEYINPUT105), .B2(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(KEYINPUT105), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n640_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n640_), .B2(new_n651_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  AND4_X1   g454(.A1(G43gat), .A2(new_n627_), .A3(new_n405_), .A4(new_n628_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G43gat), .B1(new_n634_), .B2(new_n405_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n656_), .A2(KEYINPUT47), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT47), .B1(new_n656_), .B2(new_n657_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1330gat));
  AOI21_X1  g459(.A(G50gat), .B1(new_n634_), .B2(new_n362_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n627_), .A2(new_n628_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n362_), .A2(G50gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(G1331gat));
  NAND2_X1  g463(.A1(new_n580_), .A2(new_n235_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n472_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n618_), .A2(new_n631_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n587_), .A2(KEYINPUT107), .A3(new_n666_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(G57gat), .A3(new_n393_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n618_), .A2(new_n235_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n581_), .B1(new_n676_), .B2(KEYINPUT106), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n618_), .A2(new_n678_), .A3(new_n235_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n543_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G57gat), .B1(new_n680_), .B2(new_n393_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n674_), .A2(new_n675_), .A3(new_n681_), .ZN(G1332gat));
  INV_X1    g481(.A(G64gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n683_), .A3(new_n325_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n671_), .A2(new_n325_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G64gat), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1333gat));
  INV_X1    g488(.A(G71gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n680_), .A2(new_n690_), .A3(new_n405_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n669_), .A2(new_n670_), .A3(new_n405_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT49), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G71gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G71gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n691_), .B(KEYINPUT109), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1334gat));
  NAND3_X1  g499(.A1(new_n680_), .A2(new_n353_), .A3(new_n362_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n669_), .A2(new_n670_), .A3(new_n362_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(G78gat), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G78gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n701_), .B(KEYINPUT111), .C1(new_n704_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1335gat));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n621_), .A2(new_n624_), .A3(KEYINPUT113), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT113), .B1(new_n621_), .B2(new_n624_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n665_), .A2(new_n471_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n393_), .A4(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(G85gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n392_), .A2(G85gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n631_), .A2(new_n471_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n677_), .A2(new_n719_), .A3(new_n679_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n677_), .A2(KEYINPUT112), .A3(new_n719_), .A4(new_n679_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n711_), .B1(new_n716_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n715_), .A2(G85gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n723_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT114), .B(new_n726_), .C1(new_n728_), .C2(new_n718_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1336gat));
  NAND3_X1  g529(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G92gat), .B1(new_n731_), .B2(new_n596_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n596_), .A2(G92gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n733_), .ZN(G1337gat));
  NAND4_X1  g533(.A1(new_n712_), .A2(new_n713_), .A3(new_n405_), .A4(new_n714_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(G99gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n406_), .A2(new_n487_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT51), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n735_), .A2(G99gat), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n741_), .B(new_n742_), .C1(new_n728_), .C2(new_n738_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1338gat));
  OAI211_X1 g543(.A(new_n714_), .B(new_n362_), .C1(new_n621_), .C2(new_n624_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G106gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(KEYINPUT52), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n745_), .B2(G106gat), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n361_), .A2(G106gat), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n747_), .A2(new_n749_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT53), .B1(new_n757_), .B2(new_n753_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  NAND4_X1  g558(.A1(new_n543_), .A2(new_n235_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT54), .Z(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n539_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n221_), .A2(new_n222_), .A3(new_n216_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n227_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n231_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n577_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n234_), .A2(new_n573_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n549_), .B1(new_n508_), .B2(new_n551_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n556_), .A2(KEYINPUT70), .A3(new_n550_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n547_), .A2(new_n546_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n561_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n548_), .A2(new_n558_), .A3(KEYINPUT115), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n563_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n777_), .A2(KEYINPUT116), .A3(new_n563_), .A4(new_n778_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n560_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n548_), .A2(new_n558_), .A3(KEYINPUT55), .A4(new_n559_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n781_), .A2(new_n782_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(KEYINPUT117), .B2(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n787_), .A2(new_n571_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(KEYINPUT117), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n787_), .B2(new_n571_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n571_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n788_), .B1(new_n795_), .B2(new_n789_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n770_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n769_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n770_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n787_), .A2(new_n571_), .A3(new_n790_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n784_), .A2(new_n785_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n780_), .B2(new_n779_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n572_), .B1(new_n803_), .B2(new_n782_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n804_), .B2(new_n792_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT118), .B1(new_n804_), .B2(KEYINPUT56), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n800_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT119), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n763_), .B1(new_n799_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n767_), .B1(new_n566_), .B2(new_n572_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n795_), .A2(new_n789_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n571_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT58), .B(new_n810_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n620_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n768_), .B1(new_n807_), .B2(KEYINPUT119), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n797_), .A2(new_n798_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n539_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n809_), .B(new_n817_), .C1(new_n820_), .C2(KEYINPUT57), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n761_), .B1(new_n821_), .B2(new_n472_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n363_), .A2(new_n405_), .A3(new_n393_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n234_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n823_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n799_), .A2(new_n808_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n762_), .B1(new_n829_), .B2(new_n539_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n817_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n818_), .A2(new_n819_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n763_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n471_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT59), .B(new_n828_), .C1(new_n834_), .C2(new_n761_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n827_), .A2(KEYINPUT120), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT120), .B1(new_n827_), .B2(new_n835_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n234_), .A2(G113gat), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT121), .Z(new_n840_));
  AOI21_X1  g639(.A(new_n825_), .B1(new_n838_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n827_), .A2(new_n835_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n580_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n824_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n842_), .B1(new_n581_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(KEYINPUT60), .B2(new_n842_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT122), .B1(new_n844_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n581_), .B1(new_n827_), .B2(new_n835_), .ZN(new_n851_));
  OAI221_X1 g650(.A(new_n850_), .B1(new_n845_), .B2(new_n847_), .C1(new_n851_), .C2(new_n842_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n824_), .A2(new_n854_), .A3(new_n471_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n836_), .A2(new_n837_), .A3(new_n472_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n854_), .ZN(G1342gat));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n824_), .A2(new_n858_), .A3(new_n539_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n836_), .A2(new_n837_), .A3(new_n619_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1343gat));
  NAND4_X1  g660(.A1(new_n596_), .A2(new_n406_), .A3(new_n362_), .A4(new_n393_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT123), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT124), .B1(new_n822_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n822_), .A2(KEYINPUT124), .A3(new_n863_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G141gat), .B1(new_n867_), .B2(new_n235_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n330_), .B(new_n234_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1344gat));
  OAI21_X1  g669(.A(G148gat), .B1(new_n867_), .B2(new_n581_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n331_), .B(new_n580_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1345gat));
  OAI21_X1  g672(.A(new_n471_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n867_), .B2(new_n619_), .ZN(new_n877_));
  INV_X1    g676(.A(G162gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n539_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n867_), .B2(new_n879_), .ZN(G1347gat));
  INV_X1    g679(.A(new_n822_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n325_), .A2(new_n361_), .A3(new_n407_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n234_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(new_n884_), .A3(G169gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(G169gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n882_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n234_), .A2(new_n256_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT125), .Z(new_n889_));
  OAI22_X1  g688(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n889_), .ZN(G1348gat));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n581_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n253_), .ZN(G1349gat));
  NOR2_X1   g691(.A1(new_n887_), .A2(new_n472_), .ZN(new_n893_));
  MUX2_X1   g692(.A(G183gat), .B(new_n246_), .S(new_n893_), .Z(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n887_), .B2(new_n619_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n539_), .A2(new_n247_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n887_), .B2(new_n896_), .ZN(G1351gat));
  NAND2_X1  g696(.A1(new_n430_), .A2(new_n406_), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n898_), .B(KEYINPUT126), .Z(new_n899_));
  NOR3_X1   g698(.A1(new_n822_), .A2(new_n596_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n234_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n580_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n471_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n539_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT127), .B(G218gat), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n619_), .A2(new_n911_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n900_), .B2(new_n912_), .ZN(G1355gat));
endmodule


