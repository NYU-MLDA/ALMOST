//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT84), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n213_), .B2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(new_n205_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT84), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n207_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(KEYINPUT24), .B2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT80), .B1(new_n228_), .B2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230_));
  INV_X1    g029(.A(G190gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT26), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n231_), .B2(KEYINPUT26), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n228_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT25), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT82), .B1(new_n238_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n212_), .B2(KEYINPUT25), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n229_), .A2(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT82), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n227_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n225_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n238_), .A2(new_n246_), .A3(KEYINPUT82), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n226_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT83), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n219_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(G15gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT30), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n259_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT85), .B1(new_n265_), .B2(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n264_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273_));
  INV_X1    g072(.A(G43gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT31), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT3), .Z(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT2), .Z(new_n286_));
  OAI211_X1 g085(.A(new_n280_), .B(new_n282_), .C1(new_n284_), .C2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(KEYINPUT1), .B2(new_n280_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(KEYINPUT1), .B2(new_n280_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n283_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n285_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n267_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n291_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n270_), .A3(new_n269_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n292_), .A2(new_n271_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT93), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n295_), .B2(KEYINPUT4), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n303_), .B(new_n305_), .C1(new_n302_), .C2(new_n296_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n306_), .B2(new_n299_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(G85gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT33), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(KEYINPUT94), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n307_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n311_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n306_), .B2(new_n299_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n316_), .B(KEYINPUT95), .C1(new_n306_), .C2(new_n299_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n314_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n315_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT92), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT19), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n225_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT25), .B(G183gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT26), .B(G190gat), .Z(new_n331_));
  OAI211_X1 g130(.A(new_n328_), .B(new_n226_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n206_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT90), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n206_), .B2(new_n333_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n332_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G197gat), .B(G204gat), .Z(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(KEYINPUT21), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(KEYINPUT21), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n344_), .B(new_n345_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n343_), .A2(new_n346_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT20), .B(new_n327_), .C1(new_n338_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n259_), .A2(KEYINPUT91), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT91), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n253_), .B(new_n226_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n328_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n252_), .A2(new_n253_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n218_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n352_), .B1(new_n356_), .B2(new_n347_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n349_), .B1(new_n351_), .B2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n218_), .B(new_n350_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n338_), .B2(new_n347_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n327_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND3_X1  g166(.A1(new_n358_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT91), .B1(new_n259_), .B2(new_n350_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n356_), .A2(new_n352_), .A3(new_n347_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n348_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n370_), .B1(new_n373_), .B2(new_n362_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n324_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n368_), .A2(new_n374_), .A3(KEYINPUT92), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n323_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n307_), .A2(new_n312_), .ZN(new_n379_));
  AOI211_X1 g178(.A(new_n311_), .B(new_n300_), .C1(new_n306_), .C2(new_n299_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(new_n372_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n362_), .B1(new_n383_), .B2(new_n349_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n387_));
  AND2_X1   g186(.A1(new_n332_), .A2(new_n334_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n350_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n327_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n359_), .A2(new_n361_), .A3(new_n327_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT97), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n359_), .A2(new_n361_), .A3(KEYINPUT97), .A4(new_n327_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n382_), .B(new_n386_), .C1(new_n396_), .C2(new_n385_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n378_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n401_));
  XOR2_X1   g200(.A(G22gat), .B(G50gat), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n401_), .A2(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n400_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n347_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(G228gat), .B2(G233gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n411_), .B2(new_n347_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n410_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n417_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT88), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n416_), .A2(KEYINPUT89), .A3(new_n418_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n421_), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(new_n422_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n410_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n398_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n389_), .B1(new_n351_), .B2(new_n357_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n326_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n393_), .A2(new_n394_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n367_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n368_), .A2(KEYINPUT27), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n433_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n370_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n384_), .B2(new_n367_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT98), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT27), .B1(new_n368_), .B2(new_n374_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n444_), .A2(new_n446_), .A3(new_n381_), .A4(new_n430_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n279_), .B1(new_n432_), .B2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n430_), .A2(new_n382_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n279_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT99), .B(new_n445_), .C1(new_n439_), .C2(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT100), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT98), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT98), .B1(new_n440_), .B2(new_n442_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n446_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT99), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n444_), .A2(new_n452_), .A3(new_n446_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT100), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n451_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n448_), .B1(new_n456_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT75), .B(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT76), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n476_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n476_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n479_), .B(KEYINPUT15), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n481_), .B(KEYINPUT77), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n480_), .A2(new_n482_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G113gat), .B(G141gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(G169gat), .B(G197gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n489_), .A2(new_n492_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n465_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n500_));
  NAND2_X1  g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT65), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT10), .B(G99gat), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(G106gat), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G85gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT64), .ZN(new_n512_));
  NOR2_X1   g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n510_), .B2(KEYINPUT9), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT7), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n504_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n510_), .A2(new_n513_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n518_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n525_), .B2(new_n503_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT8), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  XOR2_X1   g329(.A(G71gat), .B(G78gat), .Z(new_n531_));
  OR2_X1    g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT67), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n500_), .B1(new_n528_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT70), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n528_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n528_), .B2(new_n543_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n544_), .A2(new_n545_), .B1(new_n528_), .B2(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n540_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n528_), .B(new_n537_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(G230gat), .A3(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT5), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT13), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n554_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n476_), .B(new_n562_), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n535_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT17), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n536_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n570_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n568_), .A2(KEYINPUT17), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n528_), .A2(new_n479_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT72), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n528_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n586_), .A2(new_n484_), .B1(new_n580_), .B2(new_n579_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n582_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT36), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT73), .Z(new_n596_));
  NAND3_X1  g395(.A1(new_n589_), .A2(new_n590_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n593_), .A2(KEYINPUT36), .A3(new_n594_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n595_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT74), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n575_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(KEYINPUT37), .A3(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND4_X1   g407(.A1(new_n499_), .A2(new_n561_), .A3(new_n574_), .A4(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n382_), .A3(new_n466_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT101), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n598_), .A2(new_n603_), .A3(KEYINPUT102), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT102), .B1(new_n598_), .B2(new_n603_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n465_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n559_), .A2(new_n560_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n574_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n620_), .A2(new_n498_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n381_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n613_), .A2(new_n614_), .A3(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(new_n462_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n467_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT39), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n609_), .A2(new_n467_), .A3(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  AOI21_X1  g432(.A(new_n261_), .B1(new_n623_), .B2(new_n279_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT41), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n609_), .A2(new_n261_), .A3(new_n279_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n623_), .B2(new_n430_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT42), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n609_), .A2(new_n638_), .A3(new_n430_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT104), .ZN(G1327gat));
  NOR3_X1   g442(.A1(new_n620_), .A2(new_n498_), .A3(new_n574_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT105), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n465_), .A2(new_n608_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n432_), .A2(new_n447_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n279_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n463_), .B1(new_n462_), .B2(new_n451_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT100), .B(new_n450_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n648_), .B1(new_n654_), .B2(new_n607_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n644_), .B1(new_n647_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n654_), .B(new_n607_), .C1(KEYINPUT105), .C2(new_n645_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n648_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n465_), .B2(new_n608_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n644_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664_), .B2(new_n381_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n617_), .A2(new_n620_), .A3(new_n574_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(new_n499_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n668_), .A2(G29gat), .A3(new_n381_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n627_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT108), .B1(new_n668_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n667_), .A2(new_n674_), .A3(new_n671_), .A4(new_n627_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n658_), .A2(new_n679_), .A3(new_n663_), .A4(new_n627_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n658_), .A2(new_n627_), .A3(new_n663_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT106), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  AND4_X1   g483(.A1(new_n678_), .A2(new_n683_), .A3(G36gat), .A4(new_n680_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n677_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n677_), .B(new_n687_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  OAI21_X1  g490(.A(new_n274_), .B1(new_n668_), .B2(new_n650_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n279_), .A2(G43gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n664_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g494(.A1(new_n668_), .A2(G50gat), .A3(new_n431_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n658_), .A2(new_n430_), .A3(new_n663_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G50gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G50gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(G1331gat));
  NOR2_X1   g500(.A1(new_n465_), .A2(new_n497_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n702_), .A2(new_n620_), .A3(new_n574_), .A4(new_n608_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT111), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n382_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n498_), .A2(new_n574_), .ZN(new_n707_));
  NOR4_X1   g506(.A1(new_n618_), .A2(new_n465_), .A3(new_n561_), .A4(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n381_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1332gat));
  NOR2_X1   g510(.A1(new_n462_), .A2(G64gat), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT112), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n704_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G64gat), .B1(new_n709_), .B2(new_n462_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT48), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT48), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n716_), .B2(new_n717_), .ZN(G1333gat));
  INV_X1    g517(.A(G71gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n708_), .B2(new_n279_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT49), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n279_), .A2(new_n719_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT113), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n704_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n708_), .B2(new_n430_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n704_), .A2(new_n726_), .A3(new_n430_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1335gat));
  NAND2_X1  g529(.A1(new_n620_), .A2(new_n621_), .ZN(new_n731_));
  NOR4_X1   g530(.A1(new_n465_), .A2(new_n617_), .A3(new_n731_), .A4(new_n497_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT114), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n508_), .A3(new_n382_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n662_), .B(KEYINPUT115), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n497_), .A3(new_n731_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n382_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n737_), .B2(new_n508_), .ZN(G1336gat));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n509_), .A3(new_n627_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n736_), .A2(new_n627_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n509_), .ZN(G1337gat));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n279_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n650_), .A2(new_n506_), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n742_), .A2(G99gat), .B1(new_n733_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(G1338gat));
  INV_X1    g545(.A(G106gat), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n731_), .A2(new_n431_), .A3(new_n497_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n662_), .B2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT52), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n747_), .A3(new_n430_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(G1339gat));
  NAND2_X1  g553(.A1(new_n707_), .A2(KEYINPUT118), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n498_), .A2(new_n756_), .A3(new_n574_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n561_), .A2(new_n608_), .A3(new_n758_), .A4(KEYINPUT119), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n755_), .A2(new_n604_), .A3(new_n606_), .A4(new_n757_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n620_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(KEYINPUT54), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n760_), .B(new_n764_), .C1(new_n761_), .C2(new_n620_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n492_), .B1(new_n480_), .B2(new_n486_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n486_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n485_), .A2(new_n769_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n489_), .A2(new_n492_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT121), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n771_), .C1(new_n556_), .C2(new_n558_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n540_), .B1(new_n539_), .B2(new_n546_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n547_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n539_), .A2(new_n546_), .A3(KEYINPUT55), .A4(new_n540_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n553_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(KEYINPUT120), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n781_), .A2(new_n787_), .A3(KEYINPUT56), .A4(new_n553_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n498_), .A2(new_n556_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n776_), .B1(new_n786_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n767_), .B1(new_n791_), .B2(new_n618_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n789_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n553_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n783_), .B(new_n554_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n796_), .B2(KEYINPUT120), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT57), .B(new_n617_), .C1(new_n797_), .C2(new_n776_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n555_), .A2(new_n771_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT58), .B(new_n799_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n607_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n792_), .A2(new_n798_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n766_), .B1(new_n805_), .B2(new_n621_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n627_), .A2(new_n381_), .A3(new_n430_), .A4(new_n650_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(G113gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n497_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n621_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n766_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n814_), .A2(new_n815_), .A3(new_n807_), .A4(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(new_n817_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n498_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n811_), .B1(new_n821_), .B2(new_n810_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n561_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n809_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n561_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n809_), .B2(new_n574_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n819_), .A2(new_n820_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n574_), .A2(G127gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT123), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n809_), .A2(new_n833_), .A3(new_n618_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n608_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n833_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT124), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n834_), .C1(new_n835_), .C2(new_n833_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n806_), .A2(new_n279_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n841_), .A2(new_n382_), .A3(new_n430_), .A4(new_n462_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n498_), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n561_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT125), .B(G148gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1345gat));
  NOR2_X1   g646(.A1(new_n842_), .A2(new_n621_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n842_), .B2(new_n608_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n617_), .A2(G162gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n842_), .B2(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(G169gat), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n806_), .A2(new_n462_), .A3(new_n450_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n497_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n857_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n855_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n497_), .A2(new_n202_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT126), .Z(new_n862_));
  OAI22_X1  g661(.A1(new_n858_), .A2(new_n859_), .B1(new_n860_), .B2(new_n862_), .ZN(G1348gat));
  NAND2_X1  g662(.A1(new_n855_), .A2(new_n620_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g664(.A1(new_n855_), .A2(new_n574_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n329_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n212_), .B2(new_n866_), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n860_), .B2(new_n608_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n617_), .A2(new_n331_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n860_), .B2(new_n870_), .ZN(G1351gat));
  NOR3_X1   g670(.A1(new_n462_), .A2(new_n382_), .A3(new_n431_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n841_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n498_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n561_), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(G204gat), .Z(G1353gat));
  NAND3_X1  g676(.A1(new_n841_), .A2(new_n574_), .A3(new_n872_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n879_));
  AND2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n878_), .B2(new_n879_), .ZN(G1354gat));
  OAI21_X1  g681(.A(G218gat), .B1(new_n873_), .B2(new_n608_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n617_), .A2(G218gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n873_), .B2(new_n884_), .ZN(G1355gat));
endmodule


