//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT20), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT22), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(G169gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n217_), .B(new_n220_), .C1(new_n221_), .C2(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(new_n217_), .A3(KEYINPUT82), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n226_), .A2(new_n228_), .A3(KEYINPUT24), .A4(new_n223_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n227_), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT82), .B1(new_n225_), .B2(new_n217_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT83), .B1(new_n233_), .B2(new_n211_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT24), .B1(new_n226_), .B2(new_n228_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n210_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n229_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT78), .B1(new_n212_), .B2(KEYINPUT25), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(G183gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT26), .B1(new_n213_), .B2(new_n214_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT26), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT80), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT26), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n248_), .A3(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n243_), .A2(new_n244_), .A3(new_n249_), .A4(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT81), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n239_), .A2(new_n242_), .B1(KEYINPUT25), .B2(new_n212_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n224_), .B1(new_n238_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT21), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n261_));
  INV_X1    g060(.A(G197gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(G204gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n258_), .B1(new_n261_), .B2(new_n259_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G211gat), .A2(G218gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n271_), .A3(new_n268_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n268_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT93), .B1(new_n273_), .B2(new_n266_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n260_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n205_), .B1(new_n257_), .B2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n260_), .A2(new_n263_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n279_), .A2(new_n265_), .B1(new_n275_), .B2(new_n260_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n221_), .A2(new_n217_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n281_), .B(new_n223_), .C1(new_n210_), .C2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT25), .B(G183gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n233_), .A2(new_n286_), .A3(new_n211_), .A4(new_n229_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n204_), .B1(new_n278_), .B2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n280_), .B(new_n224_), .C1(new_n238_), .C2(new_n256_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n283_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n290_), .A2(KEYINPUT20), .A3(new_n204_), .A4(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n289_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n224_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n252_), .A2(new_n255_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n233_), .A2(KEYINPUT83), .A3(new_n211_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n236_), .B1(new_n235_), .B2(new_n210_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n231_), .A2(new_n232_), .A3(new_n230_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n304_), .A2(new_n305_), .B1(new_n223_), .B2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n302_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(KEYINPUT20), .B(new_n288_), .C1(new_n308_), .C2(new_n280_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n204_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n301_), .B1(new_n311_), .B2(new_n293_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n202_), .B1(new_n300_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n299_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n278_), .B2(new_n288_), .ZN(new_n315_));
  AND4_X1   g114(.A1(KEYINPUT20), .A2(new_n290_), .A3(new_n310_), .A4(new_n292_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n301_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n317_), .A3(KEYINPUT27), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n257_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n320_), .B(new_n224_), .C1(new_n238_), .C2(new_n256_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT86), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n326_), .A3(new_n323_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G71gat), .B(G99gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G15gat), .B(G43gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G127gat), .A2(G134gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G127gat), .A2(G134gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT87), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n337_), .ZN(new_n339_));
  OR2_X1    g138(.A1(G113gat), .A2(G120gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G113gat), .A2(G120gat), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n334_), .A2(new_n340_), .A3(new_n335_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n338_), .B1(new_n343_), .B2(KEYINPUT87), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT31), .ZN(new_n345_));
  INV_X1    g144(.A(new_n332_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n322_), .A2(new_n326_), .A3(new_n323_), .A4(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n333_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n345_), .B1(new_n333_), .B2(new_n347_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350_));
  INV_X1    g149(.A(G155gat), .ZN(new_n351_));
  INV_X1    g150(.A(G162gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT88), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(G155gat), .B2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(KEYINPUT90), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT2), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364_));
  OAI22_X1  g163(.A1(new_n359_), .A2(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(KEYINPUT90), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT91), .B1(new_n372_), .B2(KEYINPUT2), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT91), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n364_), .A2(new_n374_), .A3(new_n363_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n357_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n372_), .A2(new_n366_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n356_), .B2(KEYINPUT1), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT1), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n356_), .A2(KEYINPUT1), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n353_), .A2(new_n384_), .A3(new_n355_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n378_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n350_), .B(new_n344_), .C1(new_n377_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT97), .ZN(new_n389_));
  INV_X1    g188(.A(new_n357_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n368_), .A2(new_n366_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n372_), .A2(KEYINPUT2), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT90), .B(KEYINPUT3), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n391_), .B(new_n392_), .C1(new_n393_), .C2(new_n366_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n373_), .A2(new_n375_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n390_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n343_), .A3(new_n386_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n368_), .A2(new_n369_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n362_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n366_), .A2(new_n368_), .B1(new_n372_), .B2(KEYINPUT2), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n373_), .A4(new_n375_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n380_), .A2(new_n382_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n353_), .A2(new_n384_), .A3(new_n355_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n390_), .A2(new_n401_), .B1(new_n404_), .B2(new_n378_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n343_), .A2(KEYINPUT87), .ZN(new_n406_));
  INV_X1    g205(.A(new_n338_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n397_), .B(KEYINPUT4), .C1(new_n405_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n396_), .A2(new_n386_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT97), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n350_), .A4(new_n344_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n389_), .A2(new_n409_), .A3(new_n411_), .A4(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n344_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n410_), .A3(new_n397_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n415_), .A2(new_n423_), .A3(new_n417_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n348_), .A2(new_n349_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT102), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT95), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n396_), .B2(new_n386_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n434_), .B2(new_n280_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n431_), .B(new_n277_), .C1(new_n405_), .C2(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT94), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n430_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n396_), .A2(new_n433_), .A3(new_n386_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n396_), .A2(new_n444_), .A3(new_n433_), .A4(new_n386_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G22gat), .B(G50gat), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n439_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n441_), .A2(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n450_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n447_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n454_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n430_), .A4(new_n452_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n319_), .A2(new_n428_), .A3(new_n429_), .A4(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n313_), .A2(new_n461_), .A3(new_n318_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n333_), .A2(new_n347_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n345_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n427_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n333_), .A2(new_n347_), .A3(new_n345_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT102), .B1(new_n463_), .B2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n462_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n455_), .A2(new_n460_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n313_), .A2(new_n472_), .A3(new_n467_), .A4(new_n318_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT101), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n461_), .A2(new_n427_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT101), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n313_), .A4(new_n318_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n426_), .A2(KEYINPUT99), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT33), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n426_), .A2(KEYINPUT99), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n311_), .A2(new_n301_), .A3(new_n293_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n389_), .A2(new_n409_), .A3(new_n410_), .A4(new_n414_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n416_), .A2(new_n411_), .A3(new_n397_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n424_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n314_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT100), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n426_), .A2(KEYINPUT99), .A3(new_n481_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n481_), .B1(new_n426_), .B2(KEYINPUT99), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n314_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT100), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n299_), .A2(KEYINPUT32), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n315_), .A2(new_n316_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n427_), .B(new_n497_), .C1(new_n496_), .C2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n489_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n461_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n478_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n348_), .A2(new_n349_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n471_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT64), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT6), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G85gat), .B(G92gat), .Z(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT10), .B(G99gat), .Z(new_n515_));
  INV_X1    g314(.A(G106gat), .ZN(new_n516_));
  AOI22_X1  g315(.A1(KEYINPUT9), .A2(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  INV_X1    g321(.A(G99gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n516_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n525_));
  OR2_X1    g324(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT65), .Z(new_n531_));
  OAI21_X1  g330(.A(new_n514_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT8), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n534_), .B(new_n514_), .C1(new_n529_), .C2(new_n531_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n521_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n539_));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n535_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n530_), .B(KEYINPUT65), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n544_), .B(new_n528_), .C1(new_n512_), .C2(new_n511_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n534_), .B1(new_n545_), .B2(new_n514_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n520_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n538_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n547_), .A2(KEYINPUT68), .A3(KEYINPUT12), .A4(new_n548_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n555_), .A2(new_n542_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n558_), .B2(new_n552_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G176gat), .ZN(new_n562_));
  INV_X1    g361(.A(G204gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n553_), .B(new_n566_), .C1(new_n558_), .C2(new_n552_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT13), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(G50gat), .ZN(new_n571_));
  AND2_X1   g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(G29gat), .A2(G36gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT69), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(G29gat), .ZN(new_n575_));
  INV_X1    g374(.A(G36gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G29gat), .A2(G36gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(G43gat), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n574_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n571_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT69), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n578_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G43gat), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n574_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(G50gat), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT15), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G15gat), .B(G22gat), .ZN(new_n593_));
  INV_X1    g392(.A(G1gat), .ZN(new_n594_));
  INV_X1    g393(.A(G8gat), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT14), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G1gat), .B(G8gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n584_), .A2(new_n589_), .A3(KEYINPUT15), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n592_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n599_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT76), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n602_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n584_), .A2(new_n599_), .A3(new_n589_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n603_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n605_), .B2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(new_n225_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n262_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n612_), .A2(KEYINPUT77), .A3(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT77), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n607_), .A2(new_n611_), .A3(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n505_), .A2(new_n570_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n548_), .B(new_n599_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT75), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT16), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(G183gat), .ZN(new_n630_));
  INV_X1    g429(.A(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n626_), .A2(new_n627_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n626_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n624_), .A2(KEYINPUT17), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n633_), .A2(new_n634_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n592_), .A2(new_n600_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT70), .B1(new_n637_), .B2(new_n536_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT70), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n547_), .A2(new_n639_), .A3(new_n600_), .A4(new_n592_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n520_), .B(new_n590_), .C1(new_n543_), .C2(new_n546_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT34), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT35), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT71), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(G134gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(new_n352_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(KEYINPUT36), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n644_), .A2(KEYINPUT35), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n646_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n641_), .B(new_n654_), .C1(new_n637_), .C2(new_n536_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n647_), .A2(new_n652_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT72), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT73), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n651_), .B(KEYINPUT36), .Z(new_n660_));
  AND2_X1   g459(.A1(new_n640_), .A2(new_n641_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n645_), .B1(new_n661_), .B2(new_n638_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n655_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n659_), .B(new_n660_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n651_), .B(KEYINPUT36), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT73), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(KEYINPUT72), .A3(new_n652_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n658_), .A2(new_n664_), .A3(new_n667_), .A4(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT37), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT74), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n665_), .A2(KEYINPUT74), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n660_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT37), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n656_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n636_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n621_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n594_), .A3(new_n427_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT38), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n674_), .A2(new_n656_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n636_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n621_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G1gat), .B1(new_n685_), .B2(new_n467_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n681_), .A2(new_n686_), .ZN(G1324gat));
  OAI21_X1  g486(.A(G8gat), .B1(new_n685_), .B2(new_n319_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT39), .ZN(new_n689_));
  INV_X1    g488(.A(new_n319_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n679_), .A2(new_n595_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n685_), .B2(new_n504_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT41), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n678_), .A2(G15gat), .A3(new_n504_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n685_), .B2(new_n461_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n461_), .A2(G22gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n678_), .B2(new_n701_), .ZN(G1327gat));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703_));
  INV_X1    g502(.A(new_n636_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n570_), .A2(new_n620_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT44), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n500_), .A2(new_n461_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n474_), .A2(new_n477_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n504_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n471_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n670_), .A2(new_n714_), .A3(new_n676_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n708_), .B1(new_n713_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n670_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n676_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n503_), .B1(new_n478_), .B2(new_n501_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n708_), .B(new_n721_), .C1(new_n722_), .C2(new_n471_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n705_), .B(new_n707_), .C1(new_n718_), .C2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n705_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n715_), .A2(new_n716_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n505_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n728_), .B2(new_n723_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n730_));
  OAI21_X1  g529(.A(new_n725_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n427_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n703_), .B1(new_n732_), .B2(G29gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT105), .B(new_n575_), .C1(new_n731_), .C2(new_n427_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n704_), .A2(new_n682_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n621_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n427_), .A2(new_n575_), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n733_), .A2(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(G1328gat));
  NAND4_X1  g537(.A1(new_n621_), .A2(new_n576_), .A3(new_n690_), .A4(new_n735_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT45), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n741_), .B(new_n576_), .C1(new_n731_), .C2(new_n690_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n728_), .A2(new_n723_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n730_), .B1(new_n743_), .B2(new_n705_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n707_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n726_), .B(new_n745_), .C1(new_n728_), .C2(new_n723_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n690_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT106), .B1(new_n747_), .B2(G36gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n740_), .B1(new_n742_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT46), .B(new_n740_), .C1(new_n742_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1329gat));
  NOR3_X1   g552(.A1(new_n736_), .A2(G43gat), .A3(new_n504_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n731_), .A2(new_n503_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G43gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT108), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n756_), .B(new_n758_), .Z(G1330gat));
  AND2_X1   g558(.A1(new_n731_), .A2(new_n472_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n472_), .A2(new_n571_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n760_), .A2(new_n571_), .B1(new_n736_), .B2(new_n762_), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n713_), .A2(new_n620_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT110), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(new_n570_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n677_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n427_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n620_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n569_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n713_), .A2(new_n684_), .A3(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT111), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n427_), .A2(G57gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(G1332gat));
  INV_X1    g573(.A(G64gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n772_), .B2(new_n690_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT48), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n775_), .A3(new_n690_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n767_), .A2(new_n780_), .A3(new_n503_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n772_), .B2(new_n503_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(G1334gat));
  INV_X1    g584(.A(G78gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n767_), .A2(new_n786_), .A3(new_n472_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n772_), .B2(new_n472_), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n790_), .ZN(G1335gat));
  NAND3_X1  g590(.A1(new_n765_), .A2(new_n570_), .A3(new_n735_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(G85gat), .B1(new_n793_), .B2(new_n427_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n770_), .A2(new_n636_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n728_), .B2(new_n723_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n427_), .A2(G85gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n794_), .B1(new_n796_), .B2(new_n797_), .ZN(G1336gat));
  AOI21_X1  g597(.A(G92gat), .B1(new_n793_), .B2(new_n690_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n690_), .A2(G92gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n796_), .B2(new_n800_), .ZN(G1337gat));
  AOI21_X1  g600(.A(new_n523_), .B1(new_n796_), .B2(new_n503_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n515_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n504_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n802_), .B1(new_n793_), .B2(new_n804_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g605(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n461_), .B(new_n795_), .C1(new_n728_), .C2(new_n723_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n808_), .A2(KEYINPUT114), .A3(new_n516_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  INV_X1    g609(.A(new_n795_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n743_), .A2(new_n472_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n812_), .B2(G106gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT114), .B1(new_n808_), .B2(new_n516_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n810_), .A3(G106gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n472_), .A2(new_n516_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n792_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n807_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n807_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n824_), .B(new_n821_), .C1(new_n814_), .C2(new_n818_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1339gat));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n558_), .B2(new_n552_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n558_), .A2(new_n552_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n558_), .A2(new_n827_), .A3(new_n552_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n564_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT56), .B(new_n564_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n602_), .B1(new_n609_), .B2(new_n603_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n615_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n601_), .A2(new_n608_), .A3(new_n604_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n843_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n844_), .A2(new_n845_), .B1(new_n616_), .B2(new_n612_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n836_), .A2(new_n567_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n836_), .A2(KEYINPUT58), .A3(new_n567_), .A4(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n721_), .A3(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n567_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n846_), .A2(new_n568_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n682_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT57), .B(new_n682_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n851_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n636_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n677_), .A2(new_n862_), .A3(new_n569_), .A4(new_n620_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT116), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n677_), .A2(new_n569_), .A3(new_n620_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT54), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n859_), .A2(new_n868_), .A3(new_n636_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n504_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(KEYINPUT119), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(KEYINPUT119), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n872_), .A2(new_n873_), .A3(KEYINPUT59), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n867_), .A2(new_n860_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT59), .ZN(new_n878_));
  INV_X1    g677(.A(G113gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n620_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n875_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n877_), .B2(new_n620_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(KEYINPUT121), .A3(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1340gat));
  INV_X1    g686(.A(new_n877_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT122), .B(G120gat), .Z(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n569_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n569_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n870_), .A2(new_n874_), .B1(new_n877_), .B2(KEYINPUT59), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n890_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n888_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1341gat));
  AOI21_X1  g696(.A(G127gat), .B1(new_n888_), .B2(new_n704_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n704_), .A2(G127gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n893_), .B2(new_n899_), .ZN(G1342gat));
  AOI21_X1  g699(.A(G134gat), .B1(new_n888_), .B2(new_n683_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n721_), .A2(G134gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n893_), .B2(new_n902_), .ZN(G1343gat));
  AOI21_X1  g702(.A(new_n503_), .B1(new_n867_), .B2(new_n860_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n904_), .A2(new_n472_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n690_), .A2(new_n467_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n769_), .A3(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g707(.A1(new_n905_), .A2(new_n570_), .A3(new_n906_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g709(.A1(new_n905_), .A2(new_n704_), .A3(new_n906_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT123), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n911_), .B(new_n913_), .ZN(G1346gat));
  AND2_X1   g713(.A1(new_n905_), .A2(new_n906_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n727_), .A2(new_n352_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n905_), .A2(new_n683_), .A3(new_n906_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n915_), .A2(new_n916_), .B1(new_n917_), .B2(new_n352_), .ZN(G1347gat));
  NAND2_X1  g717(.A1(new_n690_), .A2(new_n428_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT124), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n472_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n870_), .A2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922_), .B2(new_n620_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n922_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n769_), .A3(new_n221_), .ZN(new_n927_));
  OAI211_X1 g726(.A(KEYINPUT62), .B(G169gat), .C1(new_n922_), .C2(new_n620_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n925_), .A2(new_n927_), .A3(new_n928_), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n926_), .B2(new_n570_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n472_), .B1(new_n867_), .B2(new_n860_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n920_), .A2(new_n217_), .A3(new_n569_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  NOR2_X1   g732(.A1(new_n920_), .A2(new_n636_), .ZN(new_n934_));
  AOI21_X1  g733(.A(G183gat), .B1(new_n931_), .B2(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n636_), .A2(new_n284_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n926_), .B2(new_n936_), .ZN(G1350gat));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n870_), .A2(new_n721_), .A3(new_n921_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n939_), .A2(G190gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n683_), .A2(new_n285_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n922_), .A2(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n938_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n939_), .A2(G190gat), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n944_), .B(KEYINPUT125), .C1(new_n922_), .C2(new_n941_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n904_), .A2(new_n475_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n947_), .A2(new_n769_), .A3(new_n690_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n690_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n951_), .A2(new_n563_), .A3(new_n570_), .ZN(new_n952_));
  OAI21_X1  g751(.A(G204gat), .B1(new_n950_), .B2(new_n569_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1353gat));
  NAND2_X1  g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n947_), .A2(new_n690_), .A3(new_n704_), .A4(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n631_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n956_), .B(new_n958_), .ZN(G1354gat));
  XNOR2_X1  g758(.A(KEYINPUT126), .B(G218gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n721_), .A2(new_n960_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(KEYINPUT127), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n947_), .A2(new_n690_), .A3(new_n683_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n960_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n951_), .A2(new_n962_), .B1(new_n963_), .B2(new_n964_), .ZN(G1355gat));
endmodule


