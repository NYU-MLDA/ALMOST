//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G226gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT20), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT91), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT23), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(new_n211_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT90), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(new_n211_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n227_), .A2(new_n214_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n219_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT87), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n207_), .B1(new_n231_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n214_), .A2(new_n228_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(KEYINPUT76), .B2(new_n227_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n220_), .A2(new_n223_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n244_), .B(new_n247_), .C1(KEYINPUT76), .C2(new_n227_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n217_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n215_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n240_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n242_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT93), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n242_), .A2(KEYINPUT93), .A3(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT18), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  NAND3_X1  g062(.A1(new_n241_), .A2(new_n252_), .A3(new_n248_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT20), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n219_), .A2(new_n230_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(new_n240_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n206_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n206_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT92), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n259_), .A2(new_n263_), .A3(new_n272_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n257_), .A2(new_n258_), .B1(new_n273_), .B2(KEYINPUT92), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n263_), .B1(new_n277_), .B2(new_n272_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n203_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(KEYINPUT99), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT99), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(new_n281_), .A3(new_n263_), .A4(new_n272_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n254_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n266_), .B2(new_n240_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n269_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n269_), .B2(new_n268_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n263_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n203_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n280_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n297_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT1), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n299_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n293_), .A2(KEYINPUT2), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n294_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n293_), .A2(KEYINPUT2), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n304_), .A2(new_n310_), .A3(new_n301_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n303_), .A2(KEYINPUT94), .A3(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G113gat), .B(G120gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n312_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n311_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(KEYINPUT4), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n317_), .A2(KEYINPUT4), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT95), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n317_), .A2(new_n321_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n279_), .A2(new_n290_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n241_), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(G78gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G106gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT86), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n318_), .A2(KEYINPUT29), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n336_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n336_), .B1(new_n349_), .B2(new_n347_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n333_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n287_), .A2(KEYINPUT32), .A3(new_n263_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n263_), .A2(KEYINPUT32), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n277_), .A2(new_n272_), .A3(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n355_), .B(new_n357_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n329_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n259_), .A2(new_n274_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n272_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n288_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n323_), .A2(KEYINPUT33), .A3(new_n327_), .A4(new_n328_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n360_), .A2(new_n363_), .A3(new_n275_), .A4(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n327_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n312_), .B(new_n315_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n317_), .A2(KEYINPUT96), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(new_n322_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n366_), .A2(KEYINPUT97), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT97), .B1(new_n366_), .B2(new_n371_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n352_), .B(new_n358_), .C1(new_n365_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(G71gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G99gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT80), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT78), .B(KEYINPUT79), .Z(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n253_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n248_), .A2(KEYINPUT30), .A3(new_n252_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT81), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n391_), .A3(new_n388_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n385_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n383_), .B(new_n384_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT31), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n391_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n395_), .B1(new_n394_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT31), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n385_), .A2(new_n392_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n397_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n398_), .B1(new_n397_), .B2(new_n403_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n316_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n403_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n401_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT82), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n397_), .A2(new_n403_), .A3(new_n398_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n315_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n354_), .A2(new_n375_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT100), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n279_), .A2(new_n290_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n279_), .B2(new_n290_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n352_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n406_), .A2(new_n411_), .A3(new_n332_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n413_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G190gat), .B(G218gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G134gat), .B(G162gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT36), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G232gat), .A2(G233gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT35), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n379_), .A3(new_n340_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT6), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n430_), .B(new_n432_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n438_));
  INV_X1    g237(.A(G85gat), .ZN(new_n439_));
  INV_X1    g238(.A(G92gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT65), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT65), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(new_n445_), .A3(new_n442_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n437_), .A2(new_n438_), .A3(new_n444_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT66), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT8), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT10), .B(G99gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n340_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n434_), .A2(new_n436_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n442_), .A2(KEYINPUT9), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n441_), .A2(KEYINPUT9), .A3(new_n442_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n447_), .A2(new_n448_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n437_), .A2(KEYINPUT66), .A3(new_n444_), .A4(new_n446_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT8), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n450_), .B(new_n456_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G29gat), .B(G36gat), .Z(new_n461_));
  XOR2_X1   g260(.A(G43gat), .B(G50gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT15), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n447_), .A2(new_n448_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT8), .A3(new_n458_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(new_n463_), .A3(new_n450_), .A4(new_n456_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n427_), .A2(new_n428_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n429_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n460_), .A2(new_n464_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n429_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n468_), .A3(new_n473_), .A4(new_n469_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n424_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n422_), .A2(KEYINPUT36), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n471_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n471_), .A2(KEYINPUT70), .A3(new_n474_), .A4(new_n476_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n475_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n419_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n486_));
  XOR2_X1   g285(.A(G71gat), .B(G78gat), .Z(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G231gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G15gat), .ZN(new_n496_));
  INV_X1    g295(.A(G22gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G15gat), .A2(G22gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G1gat), .A2(G8gat), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n498_), .A2(new_n499_), .B1(KEYINPUT14), .B2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n495_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n495_), .A2(new_n501_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n492_), .B(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G127gat), .B(G155gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(G183gat), .B(G211gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT17), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n505_), .A2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n510_), .A2(KEYINPUT17), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n505_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n467_), .A2(new_n490_), .A3(new_n450_), .A4(new_n456_), .ZN(new_n516_));
  INV_X1    g315(.A(G230gat), .ZN(new_n517_));
  INV_X1    g316(.A(G233gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT12), .ZN(new_n522_));
  INV_X1    g321(.A(new_n490_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n460_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n460_), .B2(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT68), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n521_), .B(new_n528_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n460_), .A2(new_n523_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n516_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n532_), .B(new_n519_), .C1(new_n531_), .C2(new_n530_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT5), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n527_), .A2(new_n529_), .A3(new_n533_), .A4(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(KEYINPUT13), .A3(new_n541_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OR3_X1    g345(.A1(new_n502_), .A2(new_n503_), .A3(new_n463_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n495_), .B(new_n501_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n463_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n464_), .A2(new_n504_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G169gat), .B(G197gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  AND3_X1   g357(.A1(new_n553_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT74), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n558_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n554_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n551_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n553_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT74), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n546_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT101), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n483_), .A2(new_n515_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n332_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n202_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  INV_X1    g374(.A(new_n569_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n279_), .A2(new_n290_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT100), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n279_), .A2(new_n290_), .A3(new_n414_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n406_), .A2(new_n411_), .A3(new_n332_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n352_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n576_), .B1(new_n582_), .B2(new_n413_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n515_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n475_), .B2(KEYINPUT71), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n481_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n481_), .A2(new_n585_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n544_), .A2(new_n545_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n202_), .A3(new_n573_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n574_), .B1(new_n575_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n575_), .B2(new_n592_), .ZN(G1324gat));
  INV_X1    g393(.A(G8gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n580_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n572_), .A2(new_n596_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(G8gat), .ZN(new_n600_));
  AOI211_X1 g399(.A(KEYINPUT39), .B(new_n595_), .C1(new_n572_), .C2(new_n596_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n602_), .B(new_n604_), .ZN(G1325gat));
  INV_X1    g404(.A(new_n412_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n496_), .B1(new_n572_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT41), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n591_), .A2(new_n496_), .A3(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1326gat));
  XNOR2_X1  g409(.A(new_n352_), .B(KEYINPUT103), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n497_), .B1(new_n572_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT42), .Z(new_n614_));
  NOR2_X1   g413(.A1(new_n611_), .A2(G22gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT104), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n591_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(G1327gat));
  NAND2_X1  g417(.A1(new_n481_), .A2(new_n515_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n589_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n583_), .A2(new_n620_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n621_), .A2(G29gat), .A3(new_n332_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n571_), .A2(new_n584_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n481_), .A2(new_n585_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n481_), .A2(new_n585_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT43), .B(new_n626_), .C1(new_n582_), .C2(new_n413_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT43), .ZN(new_n628_));
  INV_X1    g427(.A(new_n626_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n419_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n623_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(KEYINPUT44), .B(new_n623_), .C1(new_n627_), .C2(new_n630_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT105), .B1(new_n635_), .B2(new_n573_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n633_), .A2(KEYINPUT105), .A3(new_n573_), .A4(new_n634_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(G29gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n622_), .B1(new_n636_), .B2(new_n638_), .ZN(G1328gat));
  NOR2_X1   g438(.A1(new_n580_), .A2(G36gat), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n419_), .A2(new_n569_), .A3(new_n620_), .A4(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT45), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT45), .ZN(new_n643_));
  OAI22_X1  g442(.A1(new_n642_), .A2(new_n643_), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n633_), .A2(new_n596_), .A3(new_n634_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G36gat), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n646_), .B(new_n649_), .ZN(G1329gat));
  INV_X1    g449(.A(G43gat), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n412_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n633_), .A2(new_n634_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n621_), .B2(new_n412_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n633_), .A2(new_n655_), .A3(new_n634_), .A4(new_n652_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1330gat));
  INV_X1    g461(.A(new_n621_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G50gat), .B1(new_n663_), .B2(new_n612_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n353_), .A2(G50gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n635_), .B2(new_n665_), .ZN(G1331gat));
  AOI21_X1  g465(.A(new_n569_), .B1(new_n582_), .B2(new_n413_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n589_), .A2(new_n667_), .A3(new_n584_), .A4(new_n626_), .ZN(new_n668_));
  INV_X1    g467(.A(G57gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n573_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n546_), .A2(new_n569_), .A3(new_n515_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n419_), .A2(new_n482_), .A3(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT109), .Z(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(new_n573_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n674_), .B2(new_n669_), .ZN(G1332gat));
  NOR2_X1   g474(.A1(new_n580_), .A2(G64gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT110), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n668_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n596_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT48), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G64gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G64gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(G1333gat));
  NAND3_X1  g482(.A1(new_n668_), .A2(new_n377_), .A3(new_n606_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT49), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n673_), .A2(new_n606_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G71gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT49), .B(new_n377_), .C1(new_n673_), .C2(new_n606_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1334gat));
  NAND3_X1  g488(.A1(new_n668_), .A2(new_n338_), .A3(new_n612_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT50), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n673_), .A2(new_n612_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(G78gat), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT50), .B(new_n338_), .C1(new_n673_), .C2(new_n612_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1335gat));
  NOR2_X1   g494(.A1(new_n546_), .A2(new_n619_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n667_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n439_), .A3(new_n573_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n589_), .A2(new_n576_), .A3(new_n515_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n419_), .A2(new_n629_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT43), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n419_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(KEYINPUT111), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n699_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n573_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n698_), .B1(new_n707_), .B2(new_n439_), .ZN(G1336gat));
  AOI21_X1  g507(.A(G92gat), .B1(new_n697_), .B2(new_n596_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT112), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n580_), .A2(new_n440_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n706_), .B2(new_n711_), .ZN(G1337gat));
  AOI21_X1  g511(.A(new_n379_), .B1(new_n706_), .B2(new_n606_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n606_), .A2(new_n451_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n697_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n713_), .A2(KEYINPUT51), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT51), .B1(new_n713_), .B2(new_n716_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1338gat));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n699_), .A2(new_n352_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n340_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n627_), .A2(new_n630_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT114), .B(G106gat), .C1(new_n724_), .C2(new_n721_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(KEYINPUT52), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n720_), .B(new_n727_), .C1(new_n722_), .C2(new_n340_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n667_), .A2(new_n340_), .A3(new_n353_), .A4(new_n696_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n726_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n726_), .A2(new_n733_), .A3(new_n728_), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1339gat));
  INV_X1    g534(.A(KEYINPUT118), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n569_), .A2(G113gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT117), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n550_), .A2(new_n551_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n554_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n563_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n567_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n541_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n527_), .A2(new_n747_), .A3(new_n529_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n516_), .A2(new_n520_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n530_), .A2(KEYINPUT12), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n460_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n516_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(KEYINPUT55), .A2(new_n752_), .B1(new_n753_), .B2(new_n519_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n748_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n755_), .B2(new_n538_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n757_), .B(new_n540_), .C1(new_n748_), .C2(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n746_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT58), .B(new_n746_), .C1(new_n756_), .C2(new_n758_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n629_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT115), .B1(new_n542_), .B2(new_n745_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  AOI211_X1 g564(.A(new_n765_), .B(new_n744_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n569_), .A2(new_n541_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n481_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n763_), .B1(new_n770_), .B2(KEYINPUT57), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n542_), .A2(new_n745_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n765_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n542_), .A2(KEYINPUT115), .A3(new_n745_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n769_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT57), .A3(new_n482_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n515_), .B1(new_n771_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n590_), .B2(new_n576_), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT54), .A4(new_n569_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n778_), .A2(new_n782_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n417_), .A2(new_n332_), .A3(new_n412_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT59), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n786_));
  INV_X1    g585(.A(new_n784_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n786_), .B(new_n787_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n740_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n780_), .A2(new_n781_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n775_), .A2(new_n482_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n776_), .A3(new_n763_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n790_), .B1(new_n794_), .B2(new_n515_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n786_), .B1(new_n795_), .B2(new_n787_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n626_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n791_), .A2(new_n792_), .B1(new_n762_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n584_), .B1(new_n798_), .B2(new_n776_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT59), .B(new_n784_), .C1(new_n799_), .C2(new_n790_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(KEYINPUT116), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n739_), .B1(new_n789_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n795_), .A2(new_n787_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n569_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n736_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n796_), .A2(KEYINPUT116), .A3(new_n800_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT116), .B1(new_n796_), .B2(new_n800_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n738_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n804_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT118), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n810_), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(KEYINPUT60), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(KEYINPUT119), .B2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n803_), .B(new_n815_), .C1(KEYINPUT119), .C2(new_n813_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n546_), .B1(new_n796_), .B2(new_n800_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n812_), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n803_), .B2(new_n584_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n789_), .A2(new_n801_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n515_), .A2(KEYINPUT120), .ZN(new_n821_));
  MUX2_X1   g620(.A(KEYINPUT120), .B(new_n821_), .S(G127gat), .Z(new_n822_));
  AOI21_X1  g621(.A(new_n819_), .B1(new_n820_), .B2(new_n822_), .ZN(G1342gat));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  INV_X1    g623(.A(G134gat), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n626_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n789_), .B2(new_n801_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n783_), .A2(new_n481_), .A3(new_n784_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT121), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n832_), .A3(new_n825_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n824_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n826_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n829_), .A2(new_n832_), .A3(new_n825_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n832_), .B1(new_n829_), .B2(new_n825_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(KEYINPUT122), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n840_), .ZN(G1343gat));
  NOR3_X1   g640(.A1(new_n795_), .A2(new_n352_), .A3(new_n606_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n596_), .A2(new_n332_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n576_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n291_), .ZN(G1344gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n546_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(new_n292_), .ZN(G1345gat));
  NAND3_X1  g647(.A1(new_n842_), .A2(new_n584_), .A3(new_n843_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT123), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n842_), .A2(new_n851_), .A3(new_n584_), .A4(new_n843_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1346gat));
  INV_X1    g655(.A(G162gat), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n844_), .A2(new_n857_), .A3(new_n626_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n844_), .B2(new_n482_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT124), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n861_), .B(new_n857_), .C1(new_n844_), .C2(new_n482_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n858_), .B1(new_n860_), .B2(new_n862_), .ZN(G1347gat));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n596_), .A2(new_n332_), .A3(new_n606_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT125), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n783_), .A3(new_n611_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n576_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n868_), .B2(new_n216_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n210_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT62), .B(G169gat), .C1(new_n867_), .C2(new_n576_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(G1348gat));
  INV_X1    g671(.A(new_n867_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G176gat), .B1(new_n873_), .B2(new_n589_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n795_), .A2(new_n353_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n866_), .A2(G176gat), .A3(new_n589_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1349gat));
  NOR3_X1   g676(.A1(new_n867_), .A2(new_n222_), .A3(new_n515_), .ZN(new_n878_));
  INV_X1    g677(.A(G183gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n584_), .A3(new_n866_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n873_), .A2(new_n224_), .A3(new_n481_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n629_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(new_n884_), .A3(G190gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(G190gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(G1351gat));
  INV_X1    g686(.A(G197gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n606_), .A2(new_n352_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n783_), .A2(new_n596_), .A3(new_n332_), .A4(new_n889_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n890_), .A2(KEYINPUT127), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(KEYINPUT127), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n888_), .B(new_n576_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n890_), .B(KEYINPUT127), .ZN(new_n894_));
  AOI21_X1  g693(.A(G197gat), .B1(new_n894_), .B2(new_n569_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n589_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G204gat), .ZN(new_n898_));
  INV_X1    g697(.A(G204gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n899_), .A3(new_n589_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1353gat));
  XNOR2_X1  g700(.A(KEYINPUT63), .B(G211gat), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n515_), .B(new_n902_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n903_));
  OR2_X1    g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n894_), .B2(new_n584_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1354gat));
  INV_X1    g705(.A(G218gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n894_), .A2(new_n907_), .A3(new_n481_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n626_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(new_n909_), .ZN(G1355gat));
endmodule


