//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT6), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT65), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT7), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT8), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G85gat), .B(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n210_), .B2(new_n207_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(G85gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n203_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n208_), .A2(new_n220_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n217_), .A2(KEYINPUT66), .A3(new_n224_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(new_n232_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n235_), .B(KEYINPUT68), .ZN(new_n240_));
  INV_X1    g039(.A(new_n238_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n227_), .A2(new_n228_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT12), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n242_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n225_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n227_), .A2(new_n228_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n227_), .A2(new_n228_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(new_n245_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n253_), .B2(new_n243_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G120gat), .B(G148gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(G176gat), .B(G204gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(new_n255_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n250_), .A2(new_n262_), .A3(new_n254_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n260_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT13), .B1(new_n265_), .B2(new_n266_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT71), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n266_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT13), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n267_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT81), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(G155gat), .B2(G162gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285_));
  INV_X1    g084(.A(G141gat), .ZN(new_n286_));
  INV_X1    g085(.A(G148gat), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .A4(KEYINPUT82), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT82), .B1(new_n291_), .B2(new_n285_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT80), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT83), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n302_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n293_), .A2(KEYINPUT84), .A3(new_n299_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n299_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n289_), .A3(new_n288_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n306_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n284_), .B1(new_n305_), .B2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n295_), .B(new_n297_), .C1(G141gat), .C2(G148gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n282_), .B(KEYINPUT81), .Z(new_n315_));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n283_), .B2(KEYINPUT1), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n314_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT29), .B1(new_n313_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G197gat), .B(G204gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n322_), .A2(new_n326_), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT86), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT85), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n321_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n329_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n321_), .B2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(KEYINPUT87), .B(KEYINPUT29), .C1(new_n313_), .C2(new_n320_), .ZN(new_n340_));
  AOI211_X1 g139(.A(KEYINPUT88), .B(new_n334_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n305_), .A2(new_n312_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n284_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n320_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n338_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n329_), .A3(new_n340_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n334_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n342_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n281_), .B(new_n336_), .C1(new_n341_), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n346_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G22gat), .B(G50gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT28), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n354_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n336_), .B1(new_n341_), .B2(new_n350_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n280_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n351_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n360_), .B2(new_n351_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n358_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n348_), .A2(new_n349_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT88), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n348_), .A2(new_n342_), .A3(new_n349_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n281_), .B1(new_n368_), .B2(new_n336_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n351_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT90), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n357_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n360_), .A2(new_n361_), .A3(new_n351_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT23), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G169gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT25), .B(G183gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT26), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(G190gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n385_), .B(new_n388_), .C1(new_n389_), .C2(new_n386_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OR3_X1    g194(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n390_), .A2(new_n380_), .A3(new_n395_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n384_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n383_), .A2(KEYINPUT92), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n383_), .A2(KEYINPUT92), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n381_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n389_), .A2(new_n385_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(new_n395_), .A3(new_n380_), .A4(new_n396_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n329_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n401_), .B1(new_n400_), .B2(KEYINPUT20), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n378_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n333_), .A2(new_n398_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n337_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n378_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT18), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n417_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n400_), .A2(KEYINPUT20), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT91), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n409_), .A3(new_n402_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n428_), .B2(new_n378_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n422_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n433_));
  NAND3_X1  g232(.A1(new_n413_), .A2(new_n414_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n378_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n428_), .B2(new_n378_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n422_), .B(KEYINPUT97), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n429_), .B2(new_n422_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n431_), .A2(new_n432_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n376_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G127gat), .B(G134gat), .Z(new_n442_));
  XOR2_X1   g241(.A(G113gat), .B(G120gat), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT79), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n442_), .A2(new_n443_), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n444_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n345_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n450_), .A3(KEYINPUT4), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n447_), .B(new_n454_), .C1(new_n313_), .C2(new_n320_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n448_), .A2(new_n450_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n452_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(G85gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT0), .B(G57gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT95), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n459_), .A2(KEYINPUT95), .A3(new_n464_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n468_), .A2(KEYINPUT96), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT96), .B1(new_n468_), .B2(new_n469_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT78), .ZN(new_n475_));
  XOR2_X1   g274(.A(G71gat), .B(G99gat), .Z(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n398_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(new_n447_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G43gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT77), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT30), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT31), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n483_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n473_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n441_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n412_), .A2(new_n422_), .A3(new_n417_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n422_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n463_), .B1(new_n457_), .B2(new_n453_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n467_), .A2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n467_), .A2(new_n497_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n491_), .A2(new_n496_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n429_), .B1(new_n501_), .B2(new_n423_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n436_), .A2(KEYINPUT32), .A3(new_n422_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n468_), .A2(new_n502_), .A3(new_n503_), .A4(new_n469_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n362_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n373_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n440_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n364_), .A3(new_n375_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n486_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT98), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n486_), .B1(new_n376_), .B2(new_n505_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n510_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n488_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G29gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT74), .B(G15gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(G22gat), .ZN(new_n523_));
  INV_X1    g322(.A(G1gat), .ZN(new_n524_));
  INV_X1    g323(.A(G8gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G8gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n521_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n529_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(new_n520_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n531_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n532_), .B(new_n520_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT75), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n539_), .B(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n279_), .A2(new_n517_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n521_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n225_), .A2(new_n546_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n252_), .B2(new_n520_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(new_n547_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  OR3_X1    g356(.A1(new_n554_), .A2(KEYINPUT36), .A3(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(KEYINPUT36), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n532_), .B(new_n570_), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n245_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  OR3_X1    g379(.A1(new_n573_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n569_), .A2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n545_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n524_), .A3(new_n472_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n515_), .B1(new_n514_), .B2(new_n510_), .ZN(new_n587_));
  AND4_X1   g386(.A1(new_n515_), .A2(new_n508_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n588_));
  OAI22_X1  g387(.A1(new_n587_), .A2(new_n588_), .B1(new_n441_), .B2(new_n487_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n561_), .B(KEYINPUT99), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR4_X1   g390(.A1(new_n591_), .A2(new_n279_), .A3(new_n583_), .A4(new_n544_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n592_), .A2(new_n472_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n586_), .B1(new_n524_), .B2(new_n593_), .ZN(new_n594_));
  MUX2_X1   g393(.A(new_n586_), .B(new_n594_), .S(KEYINPUT38), .Z(G1324gat));
  NOR3_X1   g394(.A1(new_n279_), .A2(new_n583_), .A3(new_n544_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n440_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n596_), .A2(new_n590_), .A3(new_n597_), .A4(new_n589_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n598_), .A2(KEYINPUT100), .A3(G8gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT100), .B1(new_n598_), .B2(G8gat), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n585_), .A2(new_n525_), .A3(new_n597_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n602_), .A2(KEYINPUT40), .A3(new_n603_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n604_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n592_), .B2(new_n486_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT41), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n585_), .A2(new_n611_), .A3(new_n486_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n376_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n592_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT42), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n585_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(new_n583_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n561_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n545_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(G29gat), .B1(new_n625_), .B2(new_n472_), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n622_), .B(new_n544_), .C1(new_n271_), .C2(new_n277_), .ZN(new_n627_));
  AND2_X1   g426(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n628_));
  NOR2_X1   g427(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n589_), .B2(new_n569_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n569_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n517_), .A2(new_n632_), .A3(new_n628_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n627_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n627_), .B(KEYINPUT44), .C1(new_n631_), .C2(new_n633_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n472_), .A2(G29gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n626_), .B1(new_n638_), .B2(new_n639_), .ZN(G1328gat));
  NOR2_X1   g439(.A1(new_n440_), .A2(G36gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n545_), .A2(new_n623_), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n597_), .A3(new_n637_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT102), .A3(G36gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(new_n644_), .B2(G36gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI221_X1 g449(.A(new_n643_), .B1(new_n648_), .B2(KEYINPUT46), .C1(new_n645_), .C2(new_n646_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  INV_X1    g451(.A(G43gat), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n511_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n636_), .A2(new_n637_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT104), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n624_), .B2(new_n511_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n636_), .A2(new_n658_), .A3(new_n637_), .A4(new_n654_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g460(.A(G50gat), .B1(new_n625_), .B2(new_n617_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n617_), .A2(G50gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n638_), .B2(new_n663_), .ZN(G1331gat));
  NAND2_X1  g463(.A1(new_n279_), .A2(new_n584_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT105), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n589_), .A2(new_n544_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G57gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n472_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n544_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n583_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n591_), .A2(new_n278_), .A3(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(new_n472_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n669_), .B2(new_n675_), .ZN(G1332gat));
  INV_X1    g475(.A(G64gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n668_), .A2(new_n677_), .A3(new_n597_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n674_), .B2(new_n597_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT48), .Z(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(new_n680_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1333gat));
  INV_X1    g484(.A(G71gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n668_), .A2(new_n686_), .A3(new_n486_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n674_), .B2(new_n486_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT49), .Z(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1334gat));
  NOR2_X1   g489(.A1(new_n376_), .A2(G78gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT108), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n668_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n674_), .A2(new_n617_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(G78gat), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G78gat), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n693_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n693_), .A2(new_n698_), .A3(KEYINPUT109), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1335gat));
  NOR2_X1   g502(.A1(new_n631_), .A2(new_n633_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n279_), .A2(new_n583_), .A3(new_n544_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n472_), .A2(G85gat), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT110), .Z(new_n709_));
  NOR4_X1   g508(.A1(new_n667_), .A2(new_n278_), .A3(new_n561_), .A4(new_n622_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(new_n472_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n707_), .A2(new_n709_), .B1(new_n711_), .B2(G85gat), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT111), .Z(G1336gat));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n218_), .A3(new_n597_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n710_), .A2(new_n597_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(G92gat), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT112), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n707_), .B2(new_n511_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n710_), .A2(new_n222_), .A3(new_n486_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n710_), .A2(new_n203_), .A3(new_n617_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n706_), .A2(new_n617_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G106gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT52), .B(new_n203_), .C1(new_n706_), .C2(new_n617_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n722_), .B(new_n728_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1339gat));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n247_), .B(new_n246_), .C1(new_n243_), .C2(KEYINPUT12), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n251_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n251_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n734_), .A2(new_n733_), .A3(new_n251_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n260_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT117), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT56), .B(new_n260_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n537_), .A2(new_n534_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n542_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n539_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n542_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n747_), .A2(KEYINPUT58), .A3(new_n265_), .A4(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n739_), .A2(new_n740_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n265_), .A2(new_n752_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n758_), .A3(new_n569_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n741_), .A2(KEYINPUT115), .A3(new_n746_), .ZN(new_n760_));
  OR3_X1    g559(.A1(new_n739_), .A2(KEYINPUT115), .A3(new_n740_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n544_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n763_), .A2(KEYINPUT116), .B1(new_n272_), .B2(new_n752_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n760_), .A2(new_n761_), .A3(new_n765_), .A4(new_n762_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n562_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n759_), .B1(new_n767_), .B2(KEYINPUT57), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n769_), .B(new_n562_), .C1(new_n764_), .C2(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n583_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT114), .B1(new_n270_), .B2(new_n672_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n275_), .A2(new_n773_), .A3(new_n673_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n632_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT54), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n473_), .B1(new_n771_), .B2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n441_), .A2(new_n511_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT118), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n781_), .A3(new_n778_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n671_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(G113gat), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n777_), .A2(KEYINPUT59), .A3(new_n778_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n784_), .B1(new_n671_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n789_), .B2(new_n784_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n783_), .A2(new_n784_), .B1(new_n788_), .B2(new_n791_), .ZN(G1340gat));
  INV_X1    g591(.A(KEYINPUT60), .ZN(new_n793_));
  AOI21_X1  g592(.A(G120gat), .B1(new_n279_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n793_), .B2(G120gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n780_), .A2(new_n782_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n278_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n797_));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(G1341gat));
  NAND3_X1  g598(.A1(new_n780_), .A2(new_n622_), .A3(new_n782_), .ZN(new_n800_));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n583_), .A2(KEYINPUT120), .ZN(new_n802_));
  MUX2_X1   g601(.A(KEYINPUT120), .B(new_n802_), .S(G127gat), .Z(new_n803_));
  AOI22_X1  g602(.A1(new_n800_), .A2(new_n801_), .B1(new_n788_), .B2(new_n803_), .ZN(G1342gat));
  INV_X1    g603(.A(new_n590_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n780_), .A2(new_n805_), .A3(new_n782_), .ZN(new_n806_));
  INV_X1    g605(.A(G134gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n569_), .A2(G134gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT121), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n806_), .A2(new_n807_), .B1(new_n788_), .B2(new_n809_), .ZN(G1343gat));
  NAND3_X1  g609(.A1(new_n617_), .A2(new_n440_), .A3(new_n511_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n777_), .A2(new_n671_), .A3(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT122), .B(G141gat), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1344gat));
  NAND3_X1  g614(.A1(new_n777_), .A2(new_n279_), .A3(new_n812_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT123), .B(G148gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1345gat));
  NAND2_X1  g617(.A1(new_n771_), .A2(new_n776_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(new_n472_), .A3(new_n622_), .A4(new_n812_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n777_), .A2(KEYINPUT124), .A3(new_n622_), .A4(new_n812_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1346gat));
  AND2_X1   g626(.A1(new_n777_), .A2(new_n812_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G162gat), .B1(new_n828_), .B2(new_n805_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n569_), .A2(G162gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT125), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n828_), .B2(new_n831_), .ZN(G1347gat));
  NOR3_X1   g631(.A1(new_n617_), .A2(new_n487_), .A3(new_n440_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n819_), .A2(new_n671_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT22), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n393_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(G1348gat));
  AND2_X1   g640(.A1(new_n819_), .A2(new_n833_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n279_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n622_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n385_), .ZN(new_n846_));
  INV_X1    g645(.A(G183gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n845_), .ZN(G1350gat));
  NAND3_X1  g647(.A1(new_n842_), .A2(new_n805_), .A3(new_n389_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n842_), .A2(new_n569_), .ZN(new_n850_));
  INV_X1    g649(.A(G190gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1351gat));
  XNOR2_X1  g651(.A(KEYINPUT126), .B(G197gat), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(G197gat), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n376_), .A2(new_n472_), .A3(new_n440_), .A4(new_n486_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n819_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n544_), .ZN(new_n858_));
  MUX2_X1   g657(.A(new_n853_), .B(new_n855_), .S(new_n858_), .Z(G1352gat));
  INV_X1    g658(.A(new_n857_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n279_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g661(.A1(new_n857_), .A2(new_n583_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT63), .B(G211gat), .Z(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT127), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n819_), .A2(new_n622_), .A3(new_n856_), .A4(new_n864_), .ZN(new_n866_));
  OR2_X1    g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n863_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n865_), .B1(KEYINPUT127), .B2(new_n868_), .ZN(G1354gat));
  OR3_X1    g668(.A1(new_n857_), .A2(G218gat), .A3(new_n590_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G218gat), .B1(new_n857_), .B2(new_n632_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1355gat));
endmodule


