//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G155gat), .B(G162gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n205_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n202_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n212_), .A2(KEYINPUT86), .B1(new_n214_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n210_), .A2(new_n223_), .A3(new_n211_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT28), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G228gat), .A2(G233gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT88), .B(G197gat), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(G197gat), .B2(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT89), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(KEYINPUT89), .A3(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G211gat), .B(G218gat), .Z(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n229_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n241_), .B2(new_n231_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n241_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n238_), .A2(KEYINPUT21), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n237_), .A2(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n227_), .B1(new_n245_), .B2(KEYINPUT87), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n226_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n222_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n249_));
  OAI21_X1  g048(.A(G78gat), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n236_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT89), .B1(new_n230_), .B2(new_n232_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n242_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n243_), .A2(new_n244_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n212_), .A2(KEYINPUT86), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n214_), .A2(new_n220_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n224_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT29), .ZN(new_n259_));
  INV_X1    g058(.A(G78gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n255_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(G106gat), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(G106gat), .B1(new_n250_), .B2(new_n261_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G22gat), .B(G50gat), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n250_), .A2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(G106gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n270_), .B2(new_n262_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n248_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n265_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n262_), .A3(new_n267_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n247_), .A3(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G8gat), .B(G36gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT90), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT20), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT91), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n290_), .B2(new_n289_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n290_), .B2(new_n289_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n292_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(G169gat), .B2(G176gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n291_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n302_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n288_), .B1(new_n311_), .B2(new_n255_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n307_), .A2(new_n309_), .B1(new_n296_), .B2(new_n300_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n253_), .A2(new_n254_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n287_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n298_), .A2(new_n301_), .B1(new_n309_), .B2(new_n307_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n245_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n255_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n285_), .A2(new_n288_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n281_), .B1(new_n315_), .B2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n314_), .B(KEYINPUT20), .C1(new_n245_), .C2(new_n316_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n286_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n280_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n323_), .A2(new_n286_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n245_), .B2(new_n316_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n319_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n285_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n280_), .B(KEYINPUT96), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT27), .B(new_n326_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n276_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n313_), .A2(KEYINPUT30), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n313_), .A2(KEYINPUT30), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n339_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n318_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n340_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G15gat), .B(G43gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT81), .B(KEYINPUT83), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT82), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n350_), .B(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n343_), .A2(new_n347_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G127gat), .B(G134gat), .Z(new_n359_));
  XOR2_X1   g158(.A(G113gat), .B(G120gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT31), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n358_), .A2(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366_));
  INV_X1    g165(.A(new_n361_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n258_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n258_), .A2(new_n367_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n221_), .A2(new_n361_), .A3(new_n224_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT4), .A3(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n371_), .A2(new_n374_), .B1(new_n375_), .B2(new_n369_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G85gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT0), .B(G57gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  OR2_X1    g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n369_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n370_), .A3(new_n368_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n365_), .A2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n338_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT33), .A4(new_n380_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT92), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n376_), .A2(KEYINPUT92), .A3(KEYINPUT33), .A4(new_n380_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n384_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n368_), .A2(new_n369_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n380_), .B1(new_n396_), .B2(new_n374_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n375_), .A2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n370_), .B1(new_n375_), .B2(new_n398_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n395_), .A2(new_n322_), .A3(new_n401_), .A4(new_n326_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n388_), .B1(new_n393_), .B2(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n322_), .A2(new_n401_), .A3(new_n326_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n391_), .A2(new_n392_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(KEYINPUT94), .A3(new_n405_), .A4(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n280_), .A2(KEYINPUT32), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n324_), .A2(new_n325_), .A3(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n385_), .B(new_n408_), .C1(new_n334_), .C2(new_n407_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n272_), .A2(new_n275_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n385_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n337_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n387_), .B1(new_n416_), .B2(new_n365_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G29gat), .B(G36gat), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(KEYINPUT73), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(KEYINPUT73), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G43gat), .B(G50gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G1gat), .B(G8gat), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT78), .B(G1gat), .ZN(new_n430_));
  INV_X1    g229(.A(G8gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT14), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G15gat), .B(G22gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n429_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n437_), .B(new_n428_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n427_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n427_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n419_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT15), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n426_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n424_), .A3(KEYINPUT15), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n440_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n436_), .A2(new_n438_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n428_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n441_), .A3(new_n418_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n444_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G113gat), .B(G141gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G169gat), .B(G197gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  AND3_X1   g257(.A1(new_n455_), .A2(KEYINPUT80), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n455_), .B2(KEYINPUT80), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n417_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G190gat), .B(G218gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(G134gat), .B(G162gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT36), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G232gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT7), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT67), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n476_), .A2(new_n474_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT68), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n476_), .A2(new_n474_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n486_), .B(new_n487_), .C1(new_n488_), .C2(new_n474_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G85gat), .A2(G92gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n491_), .A2(new_n492_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n487_), .B1(new_n488_), .B2(new_n474_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n484_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n493_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT10), .B(G99gat), .Z(new_n501_));
  AOI21_X1  g300(.A(new_n484_), .B1(new_n269_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT9), .A4(new_n507_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n492_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n502_), .B1(new_n512_), .B2(KEYINPUT65), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT65), .ZN(new_n514_));
  AOI211_X1 g313(.A(new_n514_), .B(new_n492_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT66), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT9), .B1(new_n496_), .B2(new_n506_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n511_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n505_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n514_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .A4(new_n502_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n500_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n524_), .A2(new_n427_), .B1(new_n471_), .B2(new_n470_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n500_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n501_), .A2(new_n269_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n485_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n519_), .B2(new_n514_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n522_), .B1(new_n529_), .B2(new_n521_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n513_), .A2(KEYINPUT66), .A3(new_n515_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT74), .B1(new_n532_), .B2(new_n449_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n446_), .A2(new_n448_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT74), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n524_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n473_), .B(new_n525_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(KEYINPUT74), .A3(new_n449_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n535_), .B1(new_n524_), .B2(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n473_), .B1(new_n541_), .B2(new_n525_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n467_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n525_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n472_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n466_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT76), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n537_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(KEYINPUT37), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT77), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(KEYINPUT77), .A3(new_n537_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n467_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n554_), .A2(new_n549_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n550_), .B1(new_n555_), .B2(KEYINPUT37), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT13), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT69), .ZN(new_n564_));
  XOR2_X1   g363(.A(G71gat), .B(G78gat), .Z(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(KEYINPUT11), .B2(new_n562_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n569_), .B(new_n526_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT12), .B1(new_n524_), .B2(new_n569_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  INV_X1    g373(.A(new_n569_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n532_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n572_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n532_), .A2(new_n575_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n571_), .B1(new_n578_), .B2(new_n570_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n561_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n570_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n571_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n524_), .B2(new_n569_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n574_), .B1(new_n532_), .B2(new_n575_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n524_), .A2(KEYINPUT12), .A3(new_n569_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n561_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n580_), .A2(new_n589_), .A3(KEYINPUT70), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT70), .B1(new_n580_), .B2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n557_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT70), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n577_), .A2(new_n579_), .A3(new_n561_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n588_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n580_), .A2(new_n589_), .A3(KEYINPUT70), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT13), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n439_), .A2(new_n440_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n575_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT16), .ZN(new_n606_));
  XOR2_X1   g405(.A(G183gat), .B(G211gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT17), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n604_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n604_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n556_), .A2(new_n600_), .A3(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n463_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n385_), .A3(new_n430_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  INV_X1    g420(.A(G1gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n385_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n599_), .A2(new_n461_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n599_), .A2(KEYINPUT97), .A3(new_n461_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(new_n614_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n338_), .A2(new_n386_), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n410_), .A2(new_n411_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n365_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n554_), .A2(new_n549_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(KEYINPUT98), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n626_), .A2(new_n614_), .A3(new_n627_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n634_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n623_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n620_), .B(new_n621_), .C1(new_n622_), .C2(new_n640_), .ZN(G1324gat));
  NAND3_X1  g440(.A1(new_n617_), .A2(new_n431_), .A3(new_n337_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n628_), .A2(new_n337_), .A3(new_n635_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(G8gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n643_), .B2(G8gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1325gat));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n636_), .A2(new_n639_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n631_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n365_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n656_));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n656_), .A2(KEYINPUT99), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n617_), .A2(new_n657_), .A3(new_n631_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(new_n652_), .A3(G15gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT99), .B1(new_n656_), .B2(new_n657_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(KEYINPUT41), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n660_), .A3(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n617_), .A2(new_n665_), .A3(new_n276_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n653_), .B2(new_n276_), .ZN(new_n667_));
  XOR2_X1   g466(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n555_), .A2(new_n615_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n600_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n463_), .A2(new_n673_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n674_), .A2(G29gat), .A3(new_n623_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n626_), .A2(new_n615_), .A3(new_n627_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n632_), .B2(new_n556_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n632_), .A2(new_n677_), .A3(new_n556_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n676_), .B(KEYINPUT44), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n385_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G29gat), .B1(new_n684_), .B2(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n675_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT102), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n414_), .A2(G36gat), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n673_), .A2(new_n632_), .A3(new_n461_), .A4(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT45), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT45), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n682_), .A2(new_n337_), .A3(new_n683_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(G36gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n689_), .A2(KEYINPUT102), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n698_), .B(new_n695_), .C1(new_n696_), .C2(G36gat), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n674_), .B2(new_n365_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT103), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n682_), .A2(G43gat), .A3(new_n631_), .A4(new_n683_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n709_), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  NAND4_X1  g510(.A1(new_n682_), .A2(G50gat), .A3(new_n276_), .A4(new_n683_), .ZN(new_n712_));
  INV_X1    g511(.A(G50gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n674_), .B2(new_n411_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1331gat));
  NAND3_X1  g514(.A1(new_n592_), .A2(new_n598_), .A3(new_n462_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n416_), .A2(new_n365_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n629_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT37), .B1(new_n554_), .B2(new_n549_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n550_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n719_), .A2(new_n615_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT104), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n385_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n716_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n635_), .A2(new_n614_), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n623_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1332gat));
  OAI21_X1  g528(.A(G64gat), .B1(new_n727_), .B2(new_n414_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT48), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n414_), .A2(G64gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT105), .Z(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n727_), .B2(new_n365_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n723_), .A2(new_n738_), .A3(new_n631_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n727_), .B2(new_n411_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n276_), .A2(new_n260_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT106), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n723_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1335gat));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747_));
  INV_X1    g546(.A(new_n672_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n718_), .B2(new_n748_), .ZN(new_n749_));
  NOR4_X1   g548(.A1(new_n417_), .A2(KEYINPUT107), .A3(new_n672_), .A4(new_n716_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n503_), .A3(new_n385_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n716_), .A2(new_n614_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n719_), .A2(new_n720_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n417_), .B2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n632_), .A2(new_n677_), .A3(new_n556_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n623_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n760_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n504_), .A3(new_n337_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G92gat), .B1(new_n759_), .B2(new_n414_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n751_), .A2(new_n631_), .A3(new_n501_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G99gat), .B1(new_n759_), .B2(new_n365_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n767_), .B(new_n769_), .ZN(G1338gat));
  XNOR2_X1  g569(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n276_), .B(new_n753_), .C1(new_n679_), .C2(new_n678_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G106gat), .B1(new_n772_), .B2(KEYINPUT110), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n758_), .B2(new_n276_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n411_), .A2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT109), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n777_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n758_), .A2(new_n774_), .A3(new_n276_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n772_), .A2(KEYINPUT110), .ZN(new_n784_));
  INV_X1    g583(.A(new_n771_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(G106gat), .A4(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n776_), .A2(new_n782_), .A3(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n776_), .A2(new_n782_), .A3(new_n786_), .A4(new_n788_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1339gat));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n516_), .A2(new_n523_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n796_), .A2(new_n526_), .A3(new_n569_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n576_), .B2(new_n573_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n577_), .A2(KEYINPUT55), .B1(new_n798_), .B2(new_n571_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT55), .B(new_n584_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT56), .B(new_n561_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n570_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n582_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n587_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n807_), .A3(new_n800_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n561_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n803_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n458_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n453_), .A2(new_n441_), .A3(new_n419_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n427_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n450_), .A2(new_n452_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n419_), .B1(new_n814_), .B2(new_n441_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n453_), .A2(new_n441_), .A3(new_n418_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n418_), .B1(new_n814_), .B2(new_n441_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n458_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT113), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n816_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n589_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n795_), .B1(new_n810_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n561_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n828_), .B2(new_n802_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT58), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n556_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n461_), .A2(new_n589_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n828_), .B2(new_n802_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n816_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n822_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n836_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n633_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n633_), .B(new_n841_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n831_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n755_), .A2(new_n614_), .A3(new_n462_), .A4(new_n599_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT54), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n721_), .A2(new_n846_), .A3(new_n462_), .A4(new_n599_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n843_), .A2(new_n615_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n338_), .A2(new_n385_), .A3(new_n631_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n794_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n829_), .A2(KEYINPUT58), .B1(new_n719_), .B2(new_n720_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n795_), .B(new_n824_), .C1(new_n828_), .C2(new_n802_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n842_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n836_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n810_), .B2(new_n832_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n841_), .B1(new_n855_), .B2(new_n633_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n615_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n845_), .A2(new_n847_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n849_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(KEYINPUT115), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n860_), .A3(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n850_), .A2(new_n864_), .A3(new_n461_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G113gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n859_), .A2(new_n860_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n462_), .A2(G113gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1340gat));
  NAND3_X1  g668(.A1(new_n850_), .A2(new_n864_), .A3(new_n600_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT116), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n850_), .A2(new_n864_), .A3(new_n872_), .A4(new_n600_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(G120gat), .A3(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n599_), .A2(KEYINPUT60), .ZN(new_n875_));
  MUX2_X1   g674(.A(new_n875_), .B(KEYINPUT60), .S(G120gat), .Z(new_n876_));
  NAND3_X1  g675(.A1(new_n859_), .A2(new_n860_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n877_), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n615_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n850_), .A2(new_n864_), .A3(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n867_), .B2(new_n615_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(KEYINPUT117), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT117), .B1(new_n881_), .B2(new_n882_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1342gat));
  AND2_X1   g684(.A1(new_n850_), .A2(new_n864_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT118), .B(G134gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n755_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n859_), .A2(new_n555_), .A3(new_n860_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n886_), .A2(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1343gat));
  NOR3_X1   g690(.A1(new_n631_), .A2(new_n623_), .A3(new_n337_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n859_), .A2(new_n276_), .A3(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n462_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT119), .B(G141gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1344gat));
  NOR2_X1   g695(.A1(new_n893_), .A2(new_n599_), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g697(.A1(new_n893_), .A2(new_n615_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT61), .B(G155gat), .Z(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  OAI21_X1  g700(.A(G162gat), .B1(new_n893_), .B2(new_n755_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n633_), .A2(G162gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n893_), .B2(new_n903_), .ZN(G1347gat));
  NOR4_X1   g703(.A1(new_n414_), .A2(new_n276_), .A3(new_n365_), .A4(new_n385_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n859_), .A2(new_n461_), .A3(new_n905_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT22), .B(G169gat), .Z(new_n907_));
  OR2_X1    g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(KEYINPUT120), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n859_), .A2(new_n911_), .A3(new_n461_), .A4(new_n905_), .ZN(new_n912_));
  AND4_X1   g711(.A1(new_n909_), .A2(new_n910_), .A3(G169gat), .A4(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(G169gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n906_), .B2(KEYINPUT120), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n909_), .B1(new_n915_), .B2(new_n912_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n908_), .B1(new_n913_), .B2(new_n916_), .ZN(G1348gat));
  NAND2_X1  g716(.A1(new_n859_), .A2(new_n905_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n600_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n305_), .B1(KEYINPUT121), .B2(G183gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n859_), .A2(new_n614_), .A3(new_n905_), .A4(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n918_), .A2(new_n615_), .ZN(new_n925_));
  INV_X1    g724(.A(G183gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT121), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n922_), .B(new_n924_), .C1(new_n925_), .C2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI211_X1 g728(.A(KEYINPUT121), .B(new_n926_), .C1(new_n918_), .C2(new_n615_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n922_), .B1(new_n930_), .B2(new_n924_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n918_), .B2(new_n755_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n555_), .A2(new_n306_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n918_), .B2(new_n934_), .ZN(G1351gat));
  AND3_X1   g734(.A1(new_n413_), .A2(new_n337_), .A3(new_n365_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n859_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n462_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(G197gat), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(KEYINPUT123), .A3(G197gat), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n938_), .B2(G197gat), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT124), .B(new_n239_), .C1(new_n937_), .C2(new_n462_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n941_), .A2(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(G1352gat));
  NOR2_X1   g745(.A1(new_n937_), .A2(new_n599_), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT125), .B(G204gat), .Z(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1353gat));
  NOR2_X1   g748(.A1(new_n937_), .A2(new_n615_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT63), .B(G211gat), .Z(new_n953_));
  NOR3_X1   g752(.A1(new_n937_), .A2(new_n615_), .A3(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT126), .B1(new_n952_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n937_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n953_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n956_), .A2(new_n614_), .A3(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n958_), .B(new_n959_), .C1(new_n950_), .C2(new_n951_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n955_), .A2(new_n960_), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n956_), .B2(new_n555_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n556_), .A2(G218gat), .ZN(new_n963_));
  XOR2_X1   g762(.A(new_n963_), .B(KEYINPUT127), .Z(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n956_), .B2(new_n964_), .ZN(G1355gat));
endmodule


