//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT76), .B(G1gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(G8gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(G15gat), .B(G22gat), .Z(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT77), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT76), .A2(G1gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT76), .A2(G1gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(G8gat), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT14), .ZN(new_n210_));
  INV_X1    g009(.A(new_n205_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n206_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n206_), .B2(new_n213_), .ZN(new_n216_));
  INV_X1    g015(.A(G36gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G29gat), .ZN(new_n218_));
  INV_X1    g017(.A(G29gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G36gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT71), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT71), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n224_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n223_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n221_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n225_), .A2(new_n228_), .A3(KEYINPUT80), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT80), .B1(new_n225_), .B2(new_n228_), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n215_), .A2(new_n216_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n214_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n204_), .A2(KEYINPUT77), .A3(new_n205_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n212_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n224_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n227_), .A2(new_n226_), .A3(new_n221_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n206_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n225_), .A2(new_n228_), .A3(KEYINPUT80), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n235_), .A2(new_n239_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n231_), .A2(KEYINPUT81), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n229_), .A2(new_n230_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n240_), .A4(new_n235_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n245_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT82), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n243_), .A2(KEYINPUT82), .A3(new_n245_), .A4(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n235_), .A2(new_n240_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n255_));
  AND3_X1   g054(.A1(new_n225_), .A2(new_n228_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(new_n244_), .A3(new_n231_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G113gat), .B(G141gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(G169gat), .B(G197gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268_));
  INV_X1    g067(.A(new_n260_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n261_), .A2(new_n268_), .A3(new_n266_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT22), .B1(new_n276_), .B2(KEYINPUT87), .ZN(new_n277_));
  INV_X1    g076(.A(G176gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G169gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n277_), .B(new_n278_), .C1(KEYINPUT87), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT88), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n276_), .A2(KEYINPUT87), .A3(KEYINPUT22), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT88), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n278_), .A4(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n283_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n282_), .A2(KEYINPUT89), .A3(new_n283_), .A4(new_n286_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  MUX2_X1   g097(.A(new_n297_), .B(KEYINPUT24), .S(new_n298_), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n292_), .B(KEYINPUT23), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n305_), .A2(KEYINPUT26), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(KEYINPUT86), .B2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n299_), .B(new_n300_), .C1(new_n303_), .C2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n296_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT90), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n296_), .A2(new_n311_), .A3(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(G15gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT30), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n313_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT92), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G120gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n319_), .A2(KEYINPUT92), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(KEYINPUT92), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT31), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n318_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n318_), .A2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G43gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  OR2_X1    g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(KEYINPUT1), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n347_));
  OR2_X1    g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n345_), .A2(new_n344_), .A3(KEYINPUT1), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n342_), .B(new_n343_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  OR3_X1    g150(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n342_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT28), .ZN(new_n363_));
  XOR2_X1   g162(.A(G22gat), .B(G50gat), .Z(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  NOR2_X1   g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT94), .B(G197gat), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(G204gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n368_), .A2(KEYINPUT21), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n367_), .A2(G204gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(G197gat), .B2(G204gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n370_), .A2(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n380_));
  AND2_X1   g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT96), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n384_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n365_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT95), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n382_), .A2(new_n383_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n363_), .B(new_n364_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n388_), .B2(KEYINPUT95), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n387_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n327_), .B(new_n359_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n327_), .A2(new_n399_), .A3(new_n359_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n397_), .B(KEYINPUT98), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n400_), .B(new_n401_), .C1(new_n395_), .C2(new_n399_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G1gat), .B(G29gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  NAND3_X1  g206(.A1(new_n398_), .A2(new_n402_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT33), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n408_), .A2(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n396_), .A2(KEYINPUT4), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n411_), .A2(new_n400_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n407_), .B1(new_n412_), .B2(new_n397_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n396_), .A2(KEYINPUT100), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n396_), .A2(KEYINPUT100), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n401_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n409_), .A2(new_n410_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n313_), .A2(new_n379_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT19), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n301_), .A2(new_n304_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n299_), .A2(new_n300_), .A3(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT22), .B(G169gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n278_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n294_), .A2(new_n283_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n379_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n418_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n379_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n310_), .A2(new_n431_), .A3(new_n312_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n379_), .B2(new_n427_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n420_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  NAND3_X1  g239(.A1(new_n430_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n431_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n443_), .A2(new_n420_), .A3(new_n428_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n421_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n441_), .A2(new_n446_), .A3(KEYINPUT97), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT97), .B1(new_n441_), .B2(new_n446_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n417_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n430_), .A2(new_n436_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT101), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT101), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n430_), .A2(new_n436_), .A3(new_n453_), .A4(new_n450_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n408_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n407_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n450_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n421_), .B1(new_n418_), .B2(new_n429_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n432_), .A2(new_n421_), .A3(new_n434_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT102), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n458_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n420_), .B1(new_n443_), .B2(new_n428_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n420_), .B2(new_n435_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT102), .A3(new_n459_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n455_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n394_), .B1(new_n449_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n441_), .A2(KEYINPUT27), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n442_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT103), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(KEYINPUT103), .A3(new_n442_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n470_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n394_), .A2(new_n458_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT27), .B1(new_n441_), .B2(new_n446_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n341_), .B1(new_n469_), .B2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n475_), .A2(new_n477_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n394_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n458_), .A4(new_n340_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n275_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G230gat), .ZN(new_n484_));
  INV_X1    g283(.A(G233gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G57gat), .B(G64gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G71gat), .B(G78gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT11), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(KEYINPUT11), .ZN(new_n490_));
  INV_X1    g289(.A(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n487_), .A2(KEYINPUT11), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n489_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G85gat), .ZN(new_n495_));
  INV_X1    g294(.A(G92gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n495_), .A2(new_n496_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT64), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n501_), .B1(new_n500_), .B2(new_n498_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n499_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n503_));
  OAI221_X1 g302(.A(new_n497_), .B1(new_n498_), .B2(new_n500_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT10), .B(G99gat), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n504_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n500_), .A2(new_n497_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517_));
  INV_X1    g316(.A(G99gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n510_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n515_), .B(new_n516_), .C1(new_n509_), .C2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT65), .B1(new_n506_), .B2(new_n508_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n505_), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n519_), .A2(new_n520_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n516_), .B1(new_n529_), .B2(new_n515_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n522_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n521_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n514_), .B1(new_n534_), .B2(new_n527_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n535_), .A2(KEYINPUT66), .A3(new_n516_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n494_), .B(new_n513_), .C1(new_n532_), .C2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT67), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT66), .B1(new_n535_), .B2(new_n516_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n530_), .A2(new_n531_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n522_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n494_), .A4(new_n513_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n494_), .B1(new_n541_), .B2(new_n513_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n486_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n537_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n513_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n552_), .B2(new_n494_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n494_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT68), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n546_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G120gat), .B(G148gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT70), .ZN(new_n561_));
  XOR2_X1   g360(.A(G176gat), .B(G204gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n546_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT13), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(KEYINPUT13), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n237_), .A2(new_n238_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT34), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n551_), .A2(new_n574_), .B1(KEYINPUT35), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n551_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  INV_X1    g379(.A(new_n576_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n578_), .B(new_n579_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n580_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n579_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n584_), .B2(new_n577_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT73), .ZN(new_n587_));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(new_n585_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT75), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n582_), .A2(new_n585_), .A3(KEYINPUT75), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n582_), .A2(new_n585_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n599_), .A3(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n494_), .B(new_n605_), .Z(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(new_n254_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n254_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT78), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT16), .ZN(new_n613_));
  XOR2_X1   g412(.A(G183gat), .B(G211gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT17), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT79), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(KEYINPUT79), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI22_X1  g422(.A1(new_n619_), .A2(new_n620_), .B1(new_n623_), .B2(new_n609_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n604_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n483_), .A2(new_n572_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n203_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n458_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n479_), .A2(new_n482_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n572_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n275_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n600_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n624_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n632_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G1gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n633_), .A2(new_n634_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n635_), .A2(new_n646_), .A3(new_n647_), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n636_), .A2(new_n640_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n480_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n638_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n651_), .A2(new_n652_), .A3(G8gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n651_), .B2(G8gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n628_), .A2(new_n629_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n480_), .A2(G8gat), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n653_), .A2(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n340_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(G15gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n661_), .B2(G15gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n660_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(KEYINPUT41), .A3(new_n663_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n630_), .A2(new_n315_), .A3(new_n340_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n666_), .A2(new_n668_), .A3(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(new_n394_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(G22gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(G22gat), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n481_), .A2(G22gat), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n673_), .A2(new_n674_), .B1(new_n655_), .B2(new_n675_), .ZN(G1327gat));
  NOR2_X1   g475(.A1(new_n609_), .A2(new_n623_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n620_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n618_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n637_), .A2(new_n679_), .A3(new_n600_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n483_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n632_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n637_), .A2(new_n679_), .A3(new_n275_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n636_), .B2(new_n604_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n604_), .ZN(new_n686_));
  AOI211_X1 g485(.A(KEYINPUT43), .B(new_n686_), .C1(new_n479_), .C2(new_n482_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT44), .B(new_n683_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n458_), .A2(new_n219_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n682_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  NAND3_X1  g493(.A1(new_n690_), .A2(new_n650_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n480_), .A2(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n483_), .A2(new_n680_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT107), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n483_), .A2(new_n700_), .A3(new_n680_), .A4(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT45), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n696_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n696_), .A2(new_n703_), .A3(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1329gat));
  NAND4_X1  g507(.A1(new_n690_), .A2(G43gat), .A3(new_n340_), .A4(new_n691_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G43gat), .B1(new_n681_), .B2(new_n340_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n713_), .B(new_n715_), .ZN(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n681_), .A2(new_n717_), .A3(new_n394_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n690_), .A2(new_n394_), .A3(new_n691_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G50gat), .B1(new_n719_), .B2(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1331gat));
  INV_X1    g522(.A(new_n275_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n572_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n649_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n458_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n636_), .A2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n625_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n458_), .B1(new_n730_), .B2(KEYINPUT111), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(KEYINPUT111), .B2(new_n730_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n732_), .B2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n726_), .B2(new_n480_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n480_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n730_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n726_), .B2(new_n341_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n341_), .A2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n730_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n726_), .B2(new_n481_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n481_), .A2(G78gat), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT112), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n730_), .B2(new_n745_), .ZN(G1335gat));
  NAND2_X1  g545(.A1(new_n636_), .A2(new_n604_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT43), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n636_), .A2(new_n684_), .A3(new_n604_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(KEYINPUT113), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n725_), .A2(new_n624_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n458_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n729_), .A2(new_n624_), .A3(new_n639_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n495_), .A3(new_n632_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1336gat));
  NAND4_X1  g558(.A1(new_n750_), .A2(new_n752_), .A3(new_n650_), .A4(new_n754_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G92gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n496_), .A3(new_n650_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT114), .ZN(G1337gat));
  NAND4_X1  g563(.A1(new_n750_), .A2(new_n752_), .A3(new_n340_), .A4(new_n754_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G99gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n340_), .A3(new_n511_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g568(.A1(new_n757_), .A2(new_n510_), .A3(new_n394_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n748_), .A2(new_n749_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n753_), .A2(new_n481_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n774_), .B2(G106gat), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT52), .B(new_n510_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n770_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n770_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n625_), .A2(new_n782_), .A3(new_n275_), .A4(new_n572_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n679_), .A2(new_n572_), .A3(new_n602_), .A4(new_n603_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n784_), .B2(new_n724_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n273_), .A2(new_n274_), .A3(new_n568_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n557_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n486_), .B1(new_n790_), .B2(new_n544_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n790_), .B2(new_n547_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n548_), .A2(new_n553_), .A3(KEYINPUT55), .A4(new_n557_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n566_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n789_), .A2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n546_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n565_), .B1(new_n546_), .B2(new_n558_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n270_), .A2(new_n271_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n266_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(KEYINPUT116), .A3(new_n266_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n259_), .A2(new_n245_), .A3(new_n231_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n804_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n811_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n270_), .A2(new_n271_), .B1(new_n817_), .B2(new_n810_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT117), .B1(new_n569_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n639_), .B1(new_n801_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n788_), .B1(new_n821_), .B2(KEYINPUT118), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n814_), .B1(new_n804_), .B2(new_n813_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n569_), .A2(KEYINPUT117), .A3(new_n818_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n566_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n273_), .A2(new_n274_), .A3(new_n568_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n823_), .B(new_n824_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(KEYINPUT118), .A3(new_n600_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n787_), .B1(new_n822_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT57), .A3(new_n600_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n805_), .A2(new_n568_), .A3(new_n812_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT58), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n835_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(KEYINPUT120), .A3(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n604_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n838_), .A2(new_n604_), .A3(KEYINPUT121), .A4(new_n842_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n834_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n827_), .A2(new_n828_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n823_), .A2(new_n824_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n600_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT119), .A3(new_n788_), .A4(new_n830_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n832_), .A2(new_n847_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n786_), .B1(new_n854_), .B2(new_n624_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n650_), .A2(new_n394_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n632_), .A3(new_n340_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(KEYINPUT59), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n852_), .A2(new_n788_), .A3(new_n830_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n843_), .A2(new_n833_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n679_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n862_), .B2(new_n786_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT123), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(new_n859_), .C1(new_n862_), .C2(new_n786_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G113gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n275_), .A2(new_n868_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n858_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n855_), .A2(new_n275_), .A3(new_n857_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(G113gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n854_), .A2(new_n624_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n786_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n857_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT122), .B(new_n868_), .C1(new_n878_), .C2(new_n275_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n870_), .B1(new_n873_), .B2(new_n879_), .ZN(G1340gat));
  AND3_X1   g679(.A1(new_n858_), .A2(new_n867_), .A3(new_n637_), .ZN(new_n881_));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n572_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(KEYINPUT60), .B2(new_n882_), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n878_), .B2(new_n884_), .ZN(G1341gat));
  NAND3_X1  g684(.A1(new_n858_), .A2(new_n867_), .A3(new_n679_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G127gat), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n878_), .A2(G127gat), .A3(new_n624_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1342gat));
  NAND3_X1  g688(.A1(new_n858_), .A2(new_n867_), .A3(new_n604_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G134gat), .ZN(new_n891_));
  OR3_X1    g690(.A1(new_n878_), .A2(G134gat), .A3(new_n600_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1343gat));
  NOR4_X1   g692(.A1(new_n650_), .A2(new_n481_), .A3(new_n340_), .A4(new_n458_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n876_), .A2(new_n894_), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n895_), .A2(G141gat), .A3(new_n275_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G141gat), .B1(new_n895_), .B2(new_n275_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1344gat));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT124), .B(G148gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n637_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n900_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n895_), .B2(new_n572_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1345gat));
  XOR2_X1   g703(.A(KEYINPUT61), .B(G155gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT125), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT126), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n899_), .A2(new_n679_), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n907_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n895_), .B2(new_n624_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1346gat));
  OR3_X1    g710(.A1(new_n895_), .A2(G162gat), .A3(new_n600_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G162gat), .B1(new_n895_), .B2(new_n686_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1347gat));
  OR2_X1    g713(.A1(new_n862_), .A2(new_n786_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n341_), .A2(new_n480_), .A3(new_n632_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n916_), .A2(new_n481_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(KEYINPUT127), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(KEYINPUT127), .B1(new_n915_), .B2(new_n917_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n724_), .A2(new_n424_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n915_), .A2(new_n724_), .A3(new_n917_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n923_), .A2(new_n924_), .A3(G169gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(G169gat), .ZN(new_n926_));
  OAI22_X1  g725(.A1(new_n921_), .A2(new_n922_), .B1(new_n925_), .B2(new_n926_), .ZN(G1348gat));
  OAI21_X1  g726(.A(new_n637_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n855_), .A2(new_n394_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n916_), .A2(G176gat), .A3(new_n637_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n928_), .A2(new_n278_), .B1(new_n929_), .B2(new_n930_), .ZN(G1349gat));
  INV_X1    g730(.A(new_n920_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n918_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n624_), .A2(new_n304_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n929_), .A2(new_n679_), .A3(new_n916_), .ZN(new_n935_));
  INV_X1    g734(.A(G183gat), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n933_), .A2(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1350gat));
  AOI21_X1  g736(.A(new_n686_), .B1(new_n932_), .B2(new_n918_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n639_), .A2(new_n301_), .ZN(new_n939_));
  OAI22_X1  g738(.A1(new_n938_), .A2(new_n305_), .B1(new_n921_), .B2(new_n939_), .ZN(G1351gat));
  NOR3_X1   g739(.A1(new_n480_), .A2(new_n340_), .A3(new_n476_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n876_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943_), .B2(new_n724_), .ZN(new_n944_));
  INV_X1    g743(.A(G197gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n942_), .A2(new_n945_), .A3(new_n275_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1352gat));
  OR3_X1    g746(.A1(new_n942_), .A2(G204gat), .A3(new_n572_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G204gat), .B1(new_n942_), .B2(new_n572_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1353gat));
  XNOR2_X1  g749(.A(KEYINPUT63), .B(G211gat), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n942_), .A2(new_n624_), .A3(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n943_), .A2(new_n679_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n952_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  OR3_X1    g754(.A1(new_n942_), .A2(G218gat), .A3(new_n600_), .ZN(new_n956_));
  OAI21_X1  g755(.A(G218gat), .B1(new_n942_), .B2(new_n686_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1355gat));
endmodule


