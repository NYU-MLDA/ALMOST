//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G43gat), .ZN(new_n203_));
  INV_X1    g002(.A(G43gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G50gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G36gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G29gat), .ZN(new_n210_));
  INV_X1    g009(.A(G29gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G36gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n208_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n208_), .B2(new_n215_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT78), .B(G1gat), .ZN(new_n220_));
  INV_X1    g019(.A(G8gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G1gat), .B(G8gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n224_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT79), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n232_), .B2(new_n225_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n219_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n219_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n229_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n217_), .A2(new_n218_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n216_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n213_), .A2(new_n214_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n206_), .A2(new_n207_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n208_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n243_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n236_), .A2(new_n237_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n238_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n242_), .B1(new_n241_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G169gat), .B(G197gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n242_), .B(new_n259_), .C1(new_n255_), .C2(new_n241_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT82), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT24), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(KEYINPUT24), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT23), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT26), .B1(new_n274_), .B2(KEYINPUT81), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n275_), .C1(new_n276_), .C2(KEYINPUT81), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n268_), .A2(new_n270_), .A3(new_n272_), .A4(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n271_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n280_), .B2(new_n271_), .ZN(new_n282_));
  OAI21_X1  g081(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n266_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n282_), .B(new_n283_), .C1(KEYINPUT22), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n278_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT30), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT84), .B(G15gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT83), .B(G43gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n265_), .B1(new_n295_), .B2(KEYINPUT86), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT85), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT31), .ZN(new_n301_));
  INV_X1    g100(.A(new_n294_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n289_), .B(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n303_), .B2(KEYINPUT87), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n265_), .B(new_n301_), .C1(new_n295_), .C2(KEYINPUT86), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  INV_X1    g114(.A(G141gat), .ZN(new_n316_));
  INV_X1    g115(.A(G148gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n318_), .A2(new_n321_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  OR2_X1    g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT88), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n316_), .A2(new_n317_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n326_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n319_), .B(new_n329_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n314_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n336_), .A2(new_n338_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n336_), .A2(new_n338_), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n328_), .A2(new_n333_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n348_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  OR3_X1    g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n342_), .A2(new_n345_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n339_), .A2(new_n341_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT90), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n339_), .A2(KEYINPUT89), .A3(new_n341_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n353_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n345_), .A2(new_n356_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT94), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n334_), .A2(KEYINPUT92), .A3(new_n300_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n300_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n348_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(KEYINPUT4), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT93), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n300_), .A2(KEYINPUT4), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(new_n348_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n367_), .A2(new_n370_), .A3(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n372_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n378_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n366_), .B1(new_n385_), .B2(KEYINPUT33), .ZN(new_n386_));
  INV_X1    g185(.A(new_n384_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n387_), .A2(new_n382_), .A3(new_n377_), .A4(new_n376_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT33), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT94), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n367_), .A2(new_n370_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n383_), .B1(new_n392_), .B2(new_n373_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n374_), .A2(new_n348_), .B1(G225gat), .B2(G233gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n371_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n314_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n285_), .A3(new_n278_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT22), .B(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(G176gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n282_), .A3(new_n269_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT26), .B(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n273_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n268_), .A2(new_n270_), .A3(new_n272_), .A4(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n397_), .B(KEYINPUT20), .C1(new_n407_), .C2(new_n396_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT19), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n396_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n410_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n286_), .A2(new_n314_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(KEYINPUT20), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT18), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n395_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n386_), .A2(new_n390_), .A3(new_n391_), .A4(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n383_), .B1(new_n378_), .B2(new_n384_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n388_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n411_), .A2(new_n415_), .A3(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n408_), .A2(new_n410_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n407_), .B2(new_n396_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n413_), .B1(new_n432_), .B2(new_n414_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n427_), .B(new_n429_), .C1(new_n428_), .C2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n365_), .B1(new_n425_), .B2(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n355_), .A2(new_n357_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT27), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n422_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n420_), .B2(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n437_), .A2(new_n442_), .A3(new_n427_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n307_), .B1(new_n436_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n305_), .A2(new_n306_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n427_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n365_), .A2(new_n442_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n264_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G120gat), .B(G148gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT5), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G176gat), .B(G204gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n452_), .B(new_n453_), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n457_));
  XOR2_X1   g256(.A(G71gat), .B(G78gat), .Z(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n457_), .A2(new_n458_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(G85gat), .A2(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT7), .ZN(new_n473_));
  INV_X1    g272(.A(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n467_), .B1(new_n472_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT67), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT66), .B(new_n467_), .C1(new_n472_), .C2(new_n478_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT8), .A4(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n464_), .A2(KEYINPUT9), .A3(new_n465_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n469_), .A2(new_n471_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n475_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n492_));
  AND2_X1   g291(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n487_), .A2(KEYINPUT65), .A3(new_n490_), .A4(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n485_), .A3(new_n490_), .A4(new_n486_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n484_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n467_), .C1(new_n472_), .C2(new_n478_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT67), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n483_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n463_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  INV_X1    g307(.A(new_n477_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n466_), .B1(new_n511_), .B2(new_n486_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n482_), .B1(new_n512_), .B2(new_n502_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT8), .B1(new_n512_), .B2(KEYINPUT66), .ZN(new_n514_));
  INV_X1    g313(.A(new_n483_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n463_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n484_), .A4(new_n500_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n507_), .A2(new_n508_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n484_), .A3(new_n500_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT68), .A3(new_n463_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(new_n525_), .A3(new_n520_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT12), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(new_n463_), .C1(new_n501_), .C2(new_n506_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n522_), .B2(new_n463_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n525_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n524_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n455_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n536_));
  OAI211_X1 g335(.A(KEYINPUT70), .B(new_n524_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n535_), .A2(new_n537_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n524_), .B(new_n455_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT71), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n450_), .B(new_n538_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n534_), .ZN(new_n543_));
  AND4_X1   g342(.A1(new_n536_), .A2(new_n543_), .A3(new_n537_), .A4(new_n454_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT13), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n522_), .A2(new_n252_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n516_), .A2(new_n235_), .A3(new_n484_), .A4(new_n500_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT72), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .A4(new_n556_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n559_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT77), .B(KEYINPUT36), .Z(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n564_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  AOI211_X1 g368(.A(new_n568_), .B(new_n569_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n561_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT37), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT80), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n253_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n463_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT16), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n580_), .A2(new_n581_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n576_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n576_), .A2(new_n582_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(new_n561_), .C1(new_n567_), .C2(new_n570_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n572_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n449_), .A2(new_n548_), .A3(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n220_), .A3(new_n427_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n444_), .A2(new_n448_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n547_), .A2(new_n264_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n586_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n571_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n446_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n599_), .A3(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(new_n442_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT97), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(KEYINPUT97), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n590_), .A2(new_n221_), .A3(new_n442_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT96), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1325gat));
  OAI21_X1  g412(.A(G15gat), .B1(new_n598_), .B2(new_n307_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT41), .Z(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n590_), .A2(new_n616_), .A3(new_n445_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1326gat));
  OAI21_X1  g417(.A(G22gat), .B1(new_n598_), .B2(new_n437_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  INV_X1    g419(.A(G22gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n590_), .A2(new_n621_), .A3(new_n365_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1327gat));
  NOR3_X1   g422(.A1(new_n547_), .A2(new_n264_), .A3(new_n586_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n572_), .A2(new_n588_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n594_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT43), .B(new_n628_), .C1(new_n444_), .C2(new_n448_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n624_), .B(KEYINPUT44), .C1(new_n627_), .C2(new_n629_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n632_), .A2(new_n427_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n571_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n586_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n547_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n449_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n427_), .A2(new_n211_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT98), .Z(new_n641_));
  OAI22_X1  g440(.A1(new_n634_), .A2(new_n211_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  NAND3_X1  g441(.A1(new_n632_), .A2(new_n442_), .A3(new_n633_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n632_), .A2(KEYINPUT99), .A3(new_n442_), .A4(new_n633_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n209_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n602_), .A2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT100), .B1(new_n639_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n449_), .A2(new_n654_), .A3(new_n638_), .A4(new_n651_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT45), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n647_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(KEYINPUT45), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n649_), .A2(new_n650_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n650_), .B1(new_n649_), .B2(new_n659_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1329gat));
  NOR2_X1   g461(.A1(new_n307_), .A2(new_n204_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n632_), .A2(new_n633_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n632_), .A2(KEYINPUT102), .A3(new_n633_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n204_), .B1(new_n639_), .B2(new_n307_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT103), .Z(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT47), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n673_), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1330gat));
  NAND3_X1  g474(.A1(new_n632_), .A2(new_n365_), .A3(new_n633_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G50gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G50gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n365_), .A2(new_n202_), .ZN(new_n680_));
  OAI22_X1  g479(.A1(new_n678_), .A2(new_n679_), .B1(new_n639_), .B2(new_n680_), .ZN(G1331gat));
  NOR2_X1   g480(.A1(new_n548_), .A2(new_n263_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n594_), .A2(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n683_), .A2(new_n596_), .A3(new_n626_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n427_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n683_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n597_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT105), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n689_), .A3(new_n597_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(G57gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n427_), .B2(KEYINPUT106), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(KEYINPUT106), .B2(new_n692_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n685_), .B1(new_n691_), .B2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n696_), .A3(new_n442_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n691_), .A2(new_n442_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(G64gat), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G64gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n684_), .A2(new_n703_), .A3(new_n445_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n688_), .A2(new_n445_), .A3(new_n690_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT49), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G71gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G71gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT108), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(G78gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n684_), .A2(new_n714_), .A3(new_n365_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n691_), .A2(new_n365_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(G78gat), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT50), .B(new_n714_), .C1(new_n691_), .C2(new_n365_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1335gat));
  OR2_X1    g519(.A1(new_n627_), .A2(new_n629_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n548_), .A2(new_n263_), .A3(new_n586_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n446_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n683_), .A2(new_n637_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n491_), .A3(new_n427_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1336gat));
  NOR2_X1   g526(.A1(new_n493_), .A2(new_n494_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n723_), .A2(new_n602_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G92gat), .B1(new_n725_), .B2(new_n442_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1337gat));
  OAI21_X1  g530(.A(G99gat), .B1(new_n723_), .B2(new_n307_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n725_), .A2(new_n445_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n475_), .A3(new_n365_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n721_), .A2(new_n365_), .A3(new_n722_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G106gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746_));
  INV_X1    g545(.A(new_n518_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n507_), .A2(KEYINPUT12), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n528_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n520_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n528_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n532_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(KEYINPUT55), .A4(new_n526_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n518_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT109), .A3(new_n521_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n745_), .A2(new_n750_), .A3(new_n753_), .A4(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n454_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n454_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n263_), .A2(new_n540_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n454_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(KEYINPUT110), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n544_), .A2(new_n545_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n230_), .A2(new_n233_), .A3(new_n219_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n240_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n260_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n241_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n772_), .B2(new_n259_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n254_), .A2(new_n775_), .A3(new_n238_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n254_), .B2(new_n238_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n240_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n262_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n762_), .A2(new_n765_), .B1(new_n766_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n743_), .B1(new_n781_), .B2(new_n571_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n538_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n454_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n784_), .A2(new_n764_), .A3(KEYINPUT110), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n757_), .A2(KEYINPUT110), .A3(new_n758_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n763_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT57), .A3(new_n635_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n540_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n779_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n777_), .A2(new_n240_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n773_), .B(new_n771_), .C1(new_n793_), .C2(new_n776_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n262_), .A4(new_n540_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n784_), .B2(new_n764_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n759_), .A2(new_n761_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT114), .A3(new_n797_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n797_), .B(KEYINPUT58), .C1(new_n784_), .C2(new_n764_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n801_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n797_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n626_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n782_), .B(new_n790_), .C1(new_n804_), .C2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n596_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n589_), .A2(new_n264_), .A3(new_n542_), .A4(new_n546_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n307_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n437_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n263_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n814_), .B1(new_n810_), .B2(new_n596_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n365_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT59), .A3(new_n817_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n264_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n827_), .B2(new_n820_), .ZN(G1340gat));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n819_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n548_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT116), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n831_), .B(new_n835_), .C1(new_n832_), .C2(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n818_), .B2(new_n596_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n840_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n823_), .A2(new_n826_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT118), .B(G127gat), .Z(new_n844_));
  NOR2_X1   g643(.A1(new_n596_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n841_), .A2(new_n842_), .B1(new_n843_), .B2(new_n845_), .ZN(G1342gat));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n819_), .A2(new_n847_), .A3(new_n571_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n628_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1343gat));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n445_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n437_), .A2(new_n442_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n446_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n855_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n824_), .A2(KEYINPUT119), .A3(new_n445_), .A4(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n264_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n316_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n548_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n317_), .ZN(G1345gat));
  OAI21_X1  g662(.A(new_n586_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT120), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n866_), .B(new_n586_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n859_), .B2(new_n628_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n635_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n859_), .B2(new_n873_), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n307_), .A2(new_n427_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n442_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n824_), .A2(new_n264_), .A3(new_n365_), .A4(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(G169gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT121), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n876_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n816_), .A2(new_n263_), .A3(new_n437_), .A4(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n879_), .A2(KEYINPUT62), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT121), .B(new_n885_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n877_), .A2(new_n400_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n884_), .B2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n879_), .A2(KEYINPUT62), .A3(new_n883_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n887_), .A4(new_n886_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(G1348gat));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n825_), .B(KEYINPUT123), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n876_), .A2(new_n401_), .A3(new_n548_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n825_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n898_), .A2(new_n548_), .A3(new_n876_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(G176gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n894_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n896_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(KEYINPUT124), .C1(G176gat), .C2(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1349gat));
  NOR2_X1   g703(.A1(new_n876_), .A2(new_n596_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G183gat), .B1(new_n895_), .B2(new_n905_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n876_), .A2(new_n273_), .A3(new_n596_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n825_), .B2(new_n907_), .ZN(G1350gat));
  NAND4_X1  g707(.A1(new_n825_), .A2(new_n404_), .A3(new_n571_), .A4(new_n880_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n898_), .A2(new_n628_), .A3(new_n876_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n274_), .ZN(G1351gat));
  NAND2_X1  g710(.A1(new_n816_), .A2(new_n307_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n365_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n263_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n547_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT125), .B(G204gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1353gat));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n586_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  INV_X1    g723(.A(new_n914_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n925_), .A2(KEYINPUT126), .A3(new_n635_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(G218gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n925_), .B2(new_n635_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n626_), .A2(G218gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT127), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n927_), .A2(new_n928_), .B1(new_n914_), .B2(new_n930_), .ZN(G1355gat));
endmodule


