//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G197gat), .B(G204gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n203_), .B1(KEYINPUT21), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT89), .B1(new_n206_), .B2(G204gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n207_), .ZN(new_n208_));
  MUX2_X1   g007(.A(new_n203_), .B(new_n205_), .S(new_n208_), .Z(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI22_X1  g014(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT85), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G155gat), .ZN(new_n223_));
  INV_X1    g022(.A(G162gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(KEYINPUT1), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n222_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G141gat), .B(G148gat), .Z(new_n232_));
  AND3_X1   g031(.A1(new_n231_), .A2(KEYINPUT86), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT86), .B1(new_n231_), .B2(new_n232_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n227_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n209_), .B1(new_n235_), .B2(KEYINPUT29), .ZN(new_n236_));
  INV_X1    g035(.A(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(G228gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(G228gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n237_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n236_), .A2(new_n243_), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n209_), .B(new_n242_), .C1(new_n235_), .C2(KEYINPUT29), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n202_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT91), .ZN(new_n247_));
  INV_X1    g046(.A(new_n209_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n227_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n231_), .A2(new_n232_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n231_), .A2(KEYINPUT86), .A3(new_n232_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n249_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n248_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n242_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n236_), .A2(new_n243_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n202_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT90), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT91), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n202_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n257_), .A2(new_n258_), .A3(new_n264_), .A4(new_n259_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n247_), .A2(new_n261_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT28), .B1(new_n235_), .B2(KEYINPUT29), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n254_), .A2(new_n268_), .A3(new_n255_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G22gat), .B(G50gat), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT92), .A4(new_n259_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n273_), .A2(new_n275_), .A3(new_n246_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT92), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n260_), .A2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n266_), .A2(new_n274_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n282_), .B(KEYINPUT80), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n289_));
  INV_X1    g088(.A(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G169gat), .B(G176gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT25), .B(G183gat), .Z(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT26), .B(G190gat), .Z(new_n295_));
  OAI221_X1 g094(.A(new_n292_), .B1(new_n293_), .B2(new_n289_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(new_n283_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n282_), .A2(KEYINPUT23), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT22), .B(G169gat), .Z(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(G176gat), .ZN(new_n303_));
  OAI22_X1  g102(.A1(new_n288_), .A2(new_n296_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n281_), .B1(new_n304_), .B2(new_n248_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n306_));
  AOI21_X1  g105(.A(G176gat), .B1(new_n306_), .B2(KEYINPUT22), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G169gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT77), .B(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT78), .B(G190gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n308_), .B1(new_n288_), .B2(new_n312_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n293_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(KEYINPUT26), .ZN(new_n318_));
  OR2_X1    g117(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321_));
  INV_X1    g120(.A(G183gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n309_), .B2(new_n321_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n315_), .B1(new_n325_), .B2(KEYINPUT79), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327_));
  AOI211_X1 g126(.A(new_n327_), .B(new_n317_), .C1(new_n320_), .C2(new_n324_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n209_), .B(new_n313_), .C1(new_n326_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n305_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n313_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n248_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n300_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n303_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n292_), .B1(new_n293_), .B2(new_n289_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n294_), .A2(new_n295_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n336_), .A2(new_n337_), .B1(new_n340_), .B2(new_n287_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n281_), .B1(new_n341_), .B2(new_n209_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n332_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G8gat), .B(G36gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n333_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n333_), .B2(new_n344_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n280_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n343_), .B1(new_n335_), .B2(new_n342_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n305_), .A2(new_n329_), .A3(new_n343_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n349_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n333_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n353_), .A2(KEYINPUT99), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT99), .B1(new_n353_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n279_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT100), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G127gat), .B(G134gat), .Z(new_n365_));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n254_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n235_), .A2(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n372_), .A2(KEYINPUT95), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT4), .ZN(new_n374_));
  INV_X1    g173(.A(new_n371_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n374_), .B(new_n375_), .C1(KEYINPUT4), .C2(new_n370_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(KEYINPUT95), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n373_), .A2(new_n376_), .A3(new_n384_), .A4(new_n377_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G71gat), .ZN(new_n389_));
  INV_X1    g188(.A(G99gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n334_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G15gat), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT82), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n394_), .B(KEYINPUT30), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n367_), .B(KEYINPUT31), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT83), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT84), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n396_), .A2(new_n397_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n399_), .A2(KEYINPUT84), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n279_), .B(KEYINPUT100), .C1(new_n360_), .C2(new_n361_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n364_), .A2(new_n387_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n402_), .A2(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n266_), .A2(new_n274_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n276_), .A2(new_n278_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n350_), .A2(KEYINPUT32), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n335_), .A2(new_n342_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n355_), .B1(new_n412_), .B2(new_n343_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n333_), .A2(new_n344_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n411_), .B(new_n413_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n415_), .A2(KEYINPUT98), .B1(KEYINPUT32), .B2(new_n350_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n386_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(KEYINPUT96), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n385_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n374_), .B(new_n371_), .C1(KEYINPUT4), .C2(new_n370_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n369_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n423_), .A2(new_n382_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n385_), .A2(new_n420_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n351_), .A2(new_n352_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n421_), .A2(new_n428_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n410_), .B1(new_n418_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n353_), .A2(new_n359_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n279_), .A2(new_n386_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n407_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n406_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G43gat), .B(G50gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G36gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G29gat), .ZN(new_n440_));
  INV_X1    g239(.A(G29gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G36gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT69), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT69), .B1(new_n440_), .B2(new_n442_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT69), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n441_), .A2(G36gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n439_), .A2(G29gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT69), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n437_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G15gat), .B(G22gat), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G8gat), .ZN(new_n455_));
  INV_X1    g254(.A(G8gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n454_), .B(new_n455_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT74), .B(G1gat), .Z(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n456_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n455_), .B1(new_n464_), .B2(new_n454_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n452_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n445_), .A2(new_n451_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n455_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n459_), .A2(new_n460_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n453_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n471_), .A3(new_n461_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n462_), .A2(new_n465_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(KEYINPUT76), .A3(new_n468_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n479_));
  AND3_X1   g278(.A1(new_n445_), .A2(new_n451_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(new_n474_), .A3(new_n466_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n478_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n436_), .A2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT101), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT6), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G85gat), .ZN(new_n504_));
  INV_X1    g303(.A(G92gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(KEYINPUT9), .A3(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n507_), .A2(KEYINPUT9), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n499_), .A2(new_n503_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n390_), .A3(new_n501_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n497_), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n495_), .A2(KEYINPUT6), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n513_), .B(new_n515_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n506_), .A2(new_n507_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n512_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n512_), .A3(new_n520_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n511_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n526_));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n526_), .A2(new_n527_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n524_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n513_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI211_X1 g337(.A(KEYINPUT8), .B(new_n519_), .C1(new_n538_), .C2(new_n499_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n510_), .B1(new_n539_), .B2(new_n521_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n532_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT65), .B1(new_n540_), .B2(new_n532_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n535_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT64), .Z(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT66), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n540_), .A2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(KEYINPUT66), .B(new_n510_), .C1(new_n539_), .C2(new_n521_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n531_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n550_), .B(KEYINPUT12), .C1(new_n529_), .C2(new_n528_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n545_), .B1(new_n524_), .B2(new_n533_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n541_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n546_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n546_), .A2(new_n557_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(KEYINPUT67), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT67), .B1(new_n563_), .B2(new_n565_), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n567_), .A2(new_n568_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n493_), .B2(KEYINPUT101), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n494_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT75), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n476_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n533_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n585_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n580_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n587_), .B2(new_n580_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n548_), .A2(new_n549_), .A3(new_n482_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n548_), .A2(KEYINPUT71), .A3(new_n482_), .A4(new_n549_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  OAI22_X1  g396(.A1(new_n540_), .A2(new_n468_), .B1(KEYINPUT35), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n605_));
  INV_X1    g404(.A(new_n603_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n606_), .A3(new_n599_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n603_), .B(new_n598_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT72), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT36), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n604_), .A2(new_n618_), .A3(new_n607_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT73), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n616_), .A2(KEYINPUT73), .A3(new_n617_), .A4(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n615_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n617_), .B1(new_n619_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n590_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n576_), .A2(KEYINPUT102), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n494_), .A2(new_n628_), .A3(new_n575_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n386_), .A2(new_n463_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n633_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n616_), .A2(new_n619_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n590_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n573_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n493_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n387_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n638_), .A3(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n360_), .A2(new_n361_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n456_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n650_), .B2(KEYINPUT39), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n652_), .A3(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT104), .B1(new_n649_), .B2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n649_), .A2(KEYINPUT105), .A3(new_n654_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n651_), .A2(new_n653_), .A3(new_n655_), .A4(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n629_), .A2(new_n456_), .A3(new_n648_), .A4(new_n632_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(KEYINPUT40), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n644_), .B2(new_n407_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  OR2_X1    g464(.A1(new_n407_), .A2(G15gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n633_), .B2(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n644_), .B2(new_n279_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n279_), .A2(G22gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n633_), .B2(new_n670_), .ZN(G1327gat));
  INV_X1    g470(.A(new_n590_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n639_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n576_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n386_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n573_), .A2(new_n590_), .A3(new_n492_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n626_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n436_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n436_), .B2(new_n680_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n678_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n436_), .A2(new_n680_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT43), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n436_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n677_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  INV_X1    g491(.A(new_n689_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n684_), .B1(new_n690_), .B2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n387_), .A2(new_n441_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n676_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n439_), .B1(new_n695_), .B2(new_n648_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n648_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n494_), .A2(new_n575_), .A3(new_n673_), .A4(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT45), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n698_), .B1(new_n699_), .B2(new_n704_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n700_), .B(new_n684_), .C1(new_n690_), .C2(new_n694_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT46), .B(new_n703_), .C1(new_n706_), .C2(new_n439_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1329gat));
  NAND2_X1  g507(.A1(new_n690_), .A2(new_n694_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(G43gat), .A3(new_n404_), .A4(new_n683_), .ZN(new_n710_));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n674_), .B2(new_n407_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n710_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n675_), .B2(new_n410_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n410_), .A2(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n695_), .B2(new_n718_), .ZN(G1331gat));
  NOR2_X1   g518(.A1(new_n573_), .A2(new_n492_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n436_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n641_), .ZN(new_n722_));
  INV_X1    g521(.A(G57gat), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n387_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n628_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n386_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n724_), .B1(new_n729_), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g529(.A(G64gat), .B1(new_n722_), .B2(new_n700_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT48), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n700_), .A2(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n725_), .B2(new_n733_), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n722_), .B2(new_n407_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n407_), .A2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n725_), .B2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n722_), .B2(new_n279_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n279_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n725_), .B2(new_n743_), .ZN(G1335gat));
  NAND2_X1  g543(.A1(new_n720_), .A2(new_n590_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n387_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n721_), .A2(new_n673_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n504_), .A3(new_n386_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1336gat));
  OAI21_X1  g550(.A(G92gat), .B1(new_n747_), .B2(new_n700_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n505_), .A3(new_n648_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n747_), .B2(new_n407_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n749_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n404_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g558(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(new_n745_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n410_), .B(new_n761_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G106gat), .B1(new_n762_), .B2(KEYINPUT112), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n746_), .B2(new_n410_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n746_), .A2(new_n764_), .A3(new_n410_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n762_), .A2(KEYINPUT112), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .A4(G106gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(new_n770_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n756_), .A2(G106gat), .A3(new_n279_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n760_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n760_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n772_), .B(new_n775_), .C1(new_n766_), .C2(new_n770_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(KEYINPUT54), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n492_), .B1(new_n778_), .B2(KEYINPUT54), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n573_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n780_), .B1(new_n628_), .B2(new_n783_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n680_), .A2(new_n782_), .A3(new_n590_), .A4(new_n779_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n492_), .A2(new_n787_), .A3(new_n565_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n492_), .B2(new_n565_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n553_), .A2(new_n556_), .A3(new_n542_), .A4(new_n535_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n792_), .B2(new_n545_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(KEYINPUT116), .A3(new_n545_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n557_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n553_), .A2(new_n554_), .A3(new_n556_), .A4(KEYINPUT55), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n562_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT56), .B(new_n562_), .C1(new_n801_), .C2(new_n793_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n791_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n473_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n483_), .A2(new_n475_), .A3(new_n466_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n489_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n491_), .B(new_n807_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n640_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT57), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n562_), .B1(new_n801_), .B2(new_n793_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n802_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n565_), .A2(new_n491_), .A3(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT58), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n819_), .B(new_n816_), .C1(new_n814_), .C2(new_n802_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n680_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n807_), .A2(new_n491_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n570_), .B2(new_n566_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n815_), .B2(new_n791_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT117), .B(new_n823_), .C1(new_n826_), .C2(new_n640_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n811_), .A2(new_n822_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n590_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n786_), .A2(new_n829_), .ZN(new_n830_));
  AND4_X1   g629(.A1(new_n386_), .A2(new_n364_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n833_));
  AND2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n832_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT119), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n833_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n839_), .B(new_n840_), .C1(new_n832_), .C2(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n492_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n832_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n846_), .B2(new_n842_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n849_), .B2(G120gat), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n852_));
  MUX2_X1   g651(.A(KEYINPUT120), .B(new_n850_), .S(new_n852_), .Z(new_n853_));
  NAND2_X1  g652(.A1(new_n832_), .A2(new_n853_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n834_), .A2(new_n837_), .A3(new_n573_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n851_), .ZN(G1341gat));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n590_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n838_), .A2(new_n841_), .A3(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n846_), .B2(new_n590_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(new_n680_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT121), .B(G134gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n838_), .A2(new_n841_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n846_), .B2(new_n639_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n648_), .A2(new_n279_), .A3(new_n387_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n628_), .A2(new_n783_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n779_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n628_), .A2(new_n783_), .A3(new_n780_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n804_), .A2(new_n808_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n810_), .B1(new_n874_), .B2(new_n639_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n875_), .A2(new_n823_), .B1(new_n821_), .B2(new_n680_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n672_), .B1(new_n876_), .B2(new_n811_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n407_), .B(new_n869_), .C1(new_n873_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n404_), .B1(new_n786_), .B2(new_n829_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT122), .A3(new_n869_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n492_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n574_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT123), .B(G148gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1345gat));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n883_), .B2(new_n672_), .ZN(new_n890_));
  AOI211_X1 g689(.A(KEYINPUT124), .B(new_n590_), .C1(new_n880_), .C2(new_n882_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n890_), .A2(new_n891_), .A3(new_n893_), .ZN(new_n894_));
  AND4_X1   g693(.A1(KEYINPUT122), .A2(new_n830_), .A3(new_n407_), .A4(new_n869_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT122), .B1(new_n881_), .B2(new_n869_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n672_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n883_), .A2(new_n889_), .A3(new_n672_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n892_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n894_), .A2(new_n900_), .ZN(G1346gat));
  INV_X1    g700(.A(new_n883_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G162gat), .B1(new_n902_), .B2(new_n862_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n883_), .A2(new_n224_), .A3(new_n640_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1347gat));
  NOR4_X1   g704(.A1(new_n407_), .A2(new_n700_), .A3(new_n410_), .A4(new_n386_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n830_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n908_), .A2(new_n842_), .A3(new_n302_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n290_), .B1(new_n907_), .B2(new_n492_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(KEYINPUT62), .B2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(KEYINPUT62), .B2(new_n910_), .ZN(G1348gat));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n574_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g713(.A1(new_n908_), .A2(new_n590_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n294_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n916_), .A2(KEYINPUT125), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n310_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(KEYINPUT125), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n908_), .B2(new_n862_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n639_), .A2(new_n295_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n908_), .B2(new_n922_), .ZN(G1351gat));
  NOR2_X1   g722(.A1(new_n279_), .A2(new_n386_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n881_), .A2(new_n924_), .A3(new_n648_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n842_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n206_), .ZN(G1352gat));
  AND4_X1   g726(.A1(new_n924_), .A2(new_n830_), .A3(new_n407_), .A4(new_n648_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n574_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g729(.A(KEYINPUT63), .B(G211gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n928_), .A2(new_n672_), .A3(new_n931_), .ZN(new_n932_));
  OAI22_X1  g731(.A1(new_n925_), .A2(new_n590_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT126), .ZN(G1354gat));
  NOR3_X1   g734(.A1(new_n925_), .A2(KEYINPUT127), .A3(new_n639_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(G218gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n925_), .B2(new_n639_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n680_), .A2(G218gat), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n937_), .A2(new_n938_), .B1(new_n928_), .B2(new_n939_), .ZN(G1355gat));
endmodule


