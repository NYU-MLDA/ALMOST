//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT79), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n208_), .B(new_n209_), .C1(G183gat), .C2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(new_n203_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n202_), .A2(new_n214_), .A3(new_n203_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n210_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT78), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223_));
  INV_X1    g022(.A(G183gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(KEYINPUT25), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n222_), .B(new_n225_), .C1(new_n226_), .C2(new_n223_), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n212_), .A2(new_n218_), .A3(new_n217_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n219_), .A2(new_n229_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n221_), .A2(new_n227_), .A3(new_n228_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n216_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n216_), .B2(new_n231_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT81), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G43gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(G15gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n239_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n236_), .A2(KEYINPUT81), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n245_), .A2(new_n237_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n246_), .B2(new_n243_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248_));
  XOR2_X1   g047(.A(G113gat), .B(G120gat), .Z(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G85gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT0), .B(G57gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT2), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT83), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(KEYINPUT83), .A3(new_n271_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT84), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n272_), .B(new_n269_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT84), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n268_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n266_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n263_), .B1(KEYINPUT1), .B2(new_n265_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(KEYINPUT1), .B2(new_n265_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n262_), .B(new_n250_), .C1(new_n280_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n250_), .ZN(new_n289_));
  AND4_X1   g088(.A1(new_n278_), .A2(new_n268_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n278_), .B1(new_n277_), .B2(new_n268_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n283_), .B(new_n289_), .C1(new_n292_), .C2(new_n266_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n250_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT91), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n280_), .A2(new_n284_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n289_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n288_), .B1(new_n299_), .B2(KEYINPUT4), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n287_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n261_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n286_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n262_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n304_), .B(new_n260_), .C1(new_n305_), .C2(new_n288_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(KEYINPUT95), .B(new_n261_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n256_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  XOR2_X1   g110(.A(G211gat), .B(G218gat), .Z(new_n312_));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G197gat), .B(G204gat), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n311_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n315_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n296_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G228gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G78gat), .B(G106gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT87), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n296_), .A2(new_n321_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n330_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n330_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n320_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n226_), .A2(KEYINPUT88), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n226_), .A2(KEYINPUT88), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n222_), .A3(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n212_), .A2(new_n218_), .A3(new_n217_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(new_n220_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n212_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n349_), .A2(new_n351_), .B1(new_n210_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n235_), .B2(new_n346_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT90), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n349_), .A2(new_n351_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n352_), .A2(new_n210_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n320_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n346_), .A2(KEYINPUT90), .A3(new_n353_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n358_), .A2(KEYINPUT20), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n320_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT89), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n216_), .A2(new_n231_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT80), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n216_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n320_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n367_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n345_), .B1(new_n359_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n375_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n367_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n373_), .A2(new_n320_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n357_), .B1(new_n381_), .B2(new_n354_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n382_), .A3(new_n344_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n355_), .A2(new_n358_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT20), .B1(new_n363_), .B2(new_n320_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n389_), .B2(new_n358_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n344_), .B(KEYINPUT98), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(KEYINPUT27), .A3(new_n383_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n386_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n340_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n310_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n380_), .A2(new_n382_), .A3(new_n398_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT96), .B1(new_n309_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404_));
  NOR4_X1   g203(.A1(new_n300_), .A2(new_n404_), .A3(new_n301_), .A4(new_n261_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n384_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT93), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n295_), .A2(new_n407_), .A3(new_n298_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n287_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n261_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT94), .B(new_n261_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n285_), .A2(new_n286_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n305_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n306_), .B2(new_n404_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n306_), .A2(new_n418_), .A3(new_n404_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n406_), .B(new_n417_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n400_), .A2(new_n401_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT96), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n308_), .A4(new_n307_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n403_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n340_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT97), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT97), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n428_), .A3(new_n340_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n309_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n340_), .A2(new_n394_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n427_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n256_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n397_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G190gat), .B(G218gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT69), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G134gat), .B(G162gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT36), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G29gat), .B(G36gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n441_), .A2(new_n442_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G43gat), .B(G50gat), .Z(new_n445_));
  OR3_X1    g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT15), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G85gat), .B(G92gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT7), .ZN(new_n456_));
  INV_X1    g255(.A(G99gat), .ZN(new_n457_));
  INV_X1    g256(.A(G106gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G99gat), .A3(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  AOI211_X1 g265(.A(new_n453_), .B(new_n455_), .C1(new_n461_), .C2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n460_), .A3(new_n459_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n453_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n454_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n452_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n463_), .A2(new_n465_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n459_), .A2(new_n460_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n455_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n468_), .A2(new_n469_), .A3(new_n454_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT65), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT10), .B(G99gat), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n458_), .ZN(new_n481_));
  INV_X1    g280(.A(G85gat), .ZN(new_n482_));
  INV_X1    g281(.A(G92gat), .ZN(new_n483_));
  OR3_X1    g282(.A1(new_n482_), .A2(new_n483_), .A3(KEYINPUT9), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n479_), .A2(new_n481_), .A3(new_n484_), .A4(new_n466_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n451_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  AOI211_X1 g286(.A(KEYINPUT66), .B(new_n487_), .C1(new_n471_), .C2(new_n477_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n450_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G232gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT34), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT35), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n491_), .A2(KEYINPUT35), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n487_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n448_), .ZN(new_n497_));
  AOI211_X1 g296(.A(new_n494_), .B(new_n495_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n489_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n492_), .A2(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n499_), .A2(new_n500_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n440_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n499_), .A2(new_n500_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n439_), .B(KEYINPUT36), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT72), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n435_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n514_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n496_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n496_), .A2(new_n518_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(KEYINPUT12), .B2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n515_), .B(KEYINPUT12), .C1(new_n516_), .C2(new_n517_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n523_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n521_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G230gat), .A2(G233gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n520_), .ZN(new_n531_));
  OAI211_X1 g330(.A(G230gat), .B(G233gat), .C1(new_n531_), .C2(new_n519_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n530_), .A2(new_n532_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(KEYINPUT13), .A3(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547_));
  INV_X1    g346(.A(G1gat), .ZN(new_n548_));
  INV_X1    g347(.A(G8gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G1gat), .B(G8gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n448_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n546_), .B(new_n555_), .C1(new_n449_), .C2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n448_), .B(new_n553_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n546_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G113gat), .B(G141gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT75), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT76), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n557_), .A2(new_n560_), .ZN(new_n570_));
  OAI22_X1  g369(.A1(new_n568_), .A2(new_n569_), .B1(new_n570_), .B2(new_n563_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n563_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n567_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT16), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n580_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n553_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(new_n518_), .Z(new_n586_));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n582_), .B(new_n583_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n587_), .B2(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n582_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n545_), .A2(new_n576_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n511_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n309_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  INV_X1    g396(.A(new_n545_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n508_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n509_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n504_), .B(new_n508_), .C1(new_n600_), .C2(new_n599_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n593_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n435_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(KEYINPUT99), .A3(new_n575_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n435_), .B2(new_n576_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n605_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n548_), .A3(new_n430_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n597_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT100), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT100), .ZN(new_n614_));
  OAI221_X1 g413(.A(new_n596_), .B1(new_n597_), .B2(new_n611_), .C1(new_n613_), .C2(new_n614_), .ZN(G1324gat));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n549_), .A3(new_n394_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n511_), .A2(new_n394_), .A3(new_n594_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n617_), .A2(KEYINPUT101), .A3(new_n618_), .A4(G8gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n549_), .B1(new_n621_), .B2(KEYINPUT39), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n617_), .A2(new_n622_), .B1(KEYINPUT101), .B2(new_n618_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n616_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n595_), .B2(new_n434_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT41), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n610_), .A2(new_n241_), .A3(new_n256_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1326gat));
  OAI21_X1  g428(.A(G22gat), .B1(new_n595_), .B2(new_n340_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n340_), .A2(G22gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT102), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n610_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(G1327gat));
  INV_X1    g434(.A(new_n593_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n509_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n545_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n430_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n598_), .A2(new_n575_), .A3(new_n593_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n602_), .A2(new_n603_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n435_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n431_), .B1(new_n426_), .B2(KEYINPUT97), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n256_), .B1(new_n649_), .B2(new_n429_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n648_), .B(new_n645_), .C1(new_n650_), .C2(new_n397_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n644_), .B1(new_n647_), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n643_), .B1(new_n652_), .B2(KEYINPUT103), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n644_), .C1(new_n647_), .C2(new_n651_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(KEYINPUT44), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n430_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n642_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  XNOR2_X1  g459(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n394_), .B(new_n657_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n394_), .B(KEYINPUT104), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n609_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n435_), .A2(new_n608_), .A3(new_n576_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n639_), .B(new_n665_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n641_), .A2(new_n671_), .A3(new_n665_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n663_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n661_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n673_), .B1(new_n662_), .B2(G36gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n661_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(KEYINPUT106), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n677_), .A2(new_n680_), .ZN(G1329gat));
  AND2_X1   g480(.A1(new_n256_), .A2(G43gat), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n656_), .A2(KEYINPUT108), .A3(new_n657_), .A4(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n657_), .B(new_n682_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT109), .B(G43gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n641_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n434_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n683_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT47), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n683_), .A2(new_n686_), .A3(new_n692_), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1330gat));
  INV_X1    g493(.A(new_n340_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G50gat), .B1(new_n641_), .B2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(G50gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n658_), .B2(new_n697_), .ZN(G1331gat));
  NAND4_X1  g497(.A1(new_n511_), .A2(new_n576_), .A3(new_n636_), .A4(new_n545_), .ZN(new_n699_));
  INV_X1    g498(.A(G57gat), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n309_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n435_), .A2(new_n575_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n604_), .A3(new_n545_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n309_), .B1(new_n703_), .B2(KEYINPUT110), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(KEYINPUT110), .B2(new_n703_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n701_), .B1(new_n705_), .B2(new_n700_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g506(.A(G64gat), .B1(new_n699_), .B2(new_n664_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT48), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n664_), .A2(G64gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n703_), .B2(new_n710_), .ZN(G1333gat));
  OAI21_X1  g510(.A(G71gat), .B1(new_n699_), .B2(new_n434_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT49), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n434_), .A2(G71gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n703_), .B2(new_n714_), .ZN(G1334gat));
  OAI21_X1  g514(.A(G78gat), .B1(new_n699_), .B2(new_n340_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT50), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n340_), .A2(G78gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n703_), .B2(new_n718_), .ZN(G1335gat));
  NAND2_X1  g518(.A1(new_n647_), .A2(new_n651_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n598_), .A2(new_n575_), .A3(new_n636_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n309_), .ZN(new_n724_));
  NOR4_X1   g523(.A1(new_n435_), .A2(new_n575_), .A3(new_n598_), .A4(new_n638_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n482_), .A3(new_n430_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1336gat));
  OAI21_X1  g526(.A(G92gat), .B1(new_n723_), .B2(new_n664_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n483_), .A3(new_n394_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1337gat));
  AND3_X1   g529(.A1(new_n725_), .A2(new_n256_), .A3(new_n480_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n722_), .A2(new_n256_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G99gat), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(KEYINPUT112), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n733_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n734_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(KEYINPUT113), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n736_), .A2(new_n738_), .B1(new_n740_), .B2(new_n742_), .ZN(G1338gat));
  NAND3_X1  g542(.A1(new_n725_), .A2(new_n458_), .A3(new_n695_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n722_), .A2(new_n695_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G106gat), .ZN(new_n747_));
  AOI211_X1 g546(.A(KEYINPUT52), .B(new_n458_), .C1(new_n722_), .C2(new_n695_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n749_), .B(new_n751_), .ZN(G1339gat));
  NAND3_X1  g551(.A1(new_n598_), .A2(new_n604_), .A3(new_n576_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT54), .Z(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT58), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT55), .B1(new_n528_), .B2(new_n529_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n530_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n528_), .A2(KEYINPUT55), .A3(new_n529_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n537_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n554_), .B1(new_n450_), .B2(new_n553_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT116), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(KEYINPUT116), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n559_), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n563_), .B1(new_n558_), .B2(new_n546_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n766_), .A2(new_n767_), .B1(new_n570_), .B2(new_n563_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(new_n540_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n539_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n761_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n756_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n760_), .A2(new_n537_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT56), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n775_), .A2(KEYINPUT58), .A3(new_n762_), .A4(new_n769_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n773_), .A2(new_n645_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n541_), .A2(new_n768_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n575_), .A2(new_n540_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT115), .B1(new_n760_), .B2(new_n537_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(KEYINPUT56), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n761_), .B1(new_n771_), .B2(KEYINPUT115), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT57), .B1(new_n784_), .B2(new_n510_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n774_), .A2(new_n786_), .A3(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(new_n780_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n783_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n778_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n509_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n777_), .B1(new_n785_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n593_), .B1(new_n793_), .B2(KEYINPUT117), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n795_), .B(new_n777_), .C1(new_n785_), .C2(new_n792_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n755_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT118), .ZN(new_n798_));
  INV_X1    g597(.A(new_n777_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n790_), .B2(new_n509_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT57), .B(new_n510_), .C1(new_n789_), .C2(new_n778_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n795_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n793_), .A2(KEYINPUT117), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n593_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n755_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n434_), .A2(new_n396_), .A3(new_n309_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n798_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n754_), .B1(new_n593_), .B2(new_n802_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n812_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n811_), .A2(KEYINPUT119), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT119), .B1(new_n811_), .B2(new_n813_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n810_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817_), .B2(new_n576_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n809_), .A2(G113gat), .A3(new_n576_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(new_n809_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT120), .B(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n821_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n598_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n810_), .A2(KEYINPUT121), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT121), .B1(new_n810_), .B2(new_n825_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n828_), .B2(new_n829_), .ZN(G1341gat));
  OAI21_X1  g629(.A(G127gat), .B1(new_n817_), .B2(new_n593_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n809_), .A2(G127gat), .A3(new_n593_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1342gat));
  OAI21_X1  g632(.A(G134gat), .B1(new_n817_), .B2(new_n646_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n809_), .A2(G134gat), .A3(new_n509_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1343gat));
  NAND2_X1  g635(.A1(new_n798_), .A2(new_n807_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n256_), .A2(new_n340_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n664_), .A2(new_n430_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n837_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842_), .B2(new_n576_), .ZN(new_n843_));
  INV_X1    g642(.A(G141gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n844_), .A3(new_n575_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1344gat));
  OAI21_X1  g645(.A(G148gat), .B1(new_n842_), .B2(new_n598_), .ZN(new_n847_));
  INV_X1    g646(.A(G148gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n841_), .A2(new_n848_), .A3(new_n545_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1345gat));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n842_), .B2(new_n593_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n841_), .A2(new_n636_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1346gat));
  AOI21_X1  g654(.A(G162gat), .B1(new_n841_), .B2(new_n510_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n645_), .A2(G162gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT122), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n841_), .B2(new_n858_), .ZN(G1347gat));
  NOR2_X1   g658(.A1(new_n664_), .A2(new_n430_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n340_), .A3(new_n256_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n811_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n576_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT123), .B1(new_n863_), .B2(new_n211_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(G169gat), .C1(new_n862_), .C2(new_n576_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(KEYINPUT62), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n202_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n867_), .B(new_n868_), .C1(KEYINPUT62), .C2(new_n864_), .ZN(G1348gat));
  INV_X1    g668(.A(new_n862_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G176gat), .B1(new_n870_), .B2(new_n545_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n837_), .A2(new_n695_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n860_), .A2(new_n256_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n873_), .A2(new_n203_), .A3(new_n598_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n872_), .B2(new_n874_), .ZN(G1349gat));
  AOI211_X1 g674(.A(new_n593_), .B(new_n862_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n593_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n837_), .A2(new_n695_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G183gat), .B1(new_n879_), .B2(new_n880_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n876_), .B1(new_n881_), .B2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n862_), .B2(new_n646_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n510_), .A2(new_n222_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n862_), .B2(new_n885_), .ZN(G1351gat));
  NAND4_X1  g685(.A1(new_n798_), .A2(new_n807_), .A3(new_n838_), .A4(new_n860_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n576_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(G197gat), .Z(G1352gat));
  INV_X1    g688(.A(G204gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n545_), .B1(KEYINPUT125), .B2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n892_), .B(new_n893_), .Z(G1353gat));
  NOR3_X1   g693(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n636_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n887_), .A2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1354gat));
  OAI21_X1  g699(.A(G218gat), .B1(new_n887_), .B2(new_n646_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n636_), .B1(new_n802_), .B2(new_n795_), .ZN(new_n902_));
  AOI211_X1 g701(.A(KEYINPUT118), .B(new_n754_), .C1(new_n902_), .C2(new_n804_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n806_), .B1(new_n805_), .B2(new_n755_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n509_), .A2(G218gat), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n905_), .A2(new_n838_), .A3(new_n860_), .A4(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n901_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n901_), .A2(new_n907_), .A3(KEYINPUT127), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1355gat));
endmodule


