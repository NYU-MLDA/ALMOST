//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT80), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(G197gat), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n211_));
  INV_X1    g010(.A(G197gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(G204gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT21), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n208_), .A2(new_n211_), .A3(G197gat), .A4(new_n209_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT21), .B1(new_n214_), .B2(new_n218_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n209_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n221_), .A2(new_n222_), .A3(G197gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT21), .B1(new_n212_), .B2(new_n207_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n215_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n219_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT73), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT73), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n227_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT73), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n236_), .A3(new_n228_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT23), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G183gat), .ZN(new_n243_));
  INV_X1    g042(.A(G190gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT26), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G190gat), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n241_), .A2(new_n243_), .A3(new_n245_), .A4(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n231_), .A2(new_n237_), .A3(new_n239_), .A4(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G169gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n238_), .B(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n226_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT19), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT71), .A2(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT26), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n246_), .A2(KEYINPUT71), .A3(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n241_), .A2(new_n243_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT72), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n231_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n255_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n226_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n257_), .A2(KEYINPUT20), .A3(new_n260_), .A4(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT20), .B1(new_n272_), .B2(new_n226_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n275_), .A2(KEYINPUT82), .B1(new_n226_), .B2(new_n256_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n277_), .B(KEYINPUT20), .C1(new_n272_), .C2(new_n226_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n205_), .B(new_n274_), .C1(new_n279_), .C2(new_n260_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n205_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n260_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n274_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(KEYINPUT83), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n287_), .B(new_n281_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n275_), .A2(KEYINPUT82), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n226_), .A2(new_n256_), .ZN(new_n291_));
  AND4_X1   g090(.A1(new_n260_), .A2(new_n290_), .A3(new_n278_), .A4(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT90), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT89), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n249_), .A2(new_n255_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n249_), .B2(new_n255_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n296_), .A2(new_n226_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT20), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n226_), .A2(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n295_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n303_), .A3(new_n273_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n292_), .B1(new_n259_), .B2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT27), .B(new_n280_), .C1(new_n305_), .C2(new_n205_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n289_), .A2(KEYINPUT95), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT95), .B1(new_n289_), .B2(new_n306_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(G155gat), .B2(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(KEYINPUT77), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT1), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(KEYINPUT77), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(G155gat), .A3(G162gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G141gat), .B(G148gat), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OR3_X1    g122(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325_));
  INV_X1    g124(.A(G141gat), .ZN(new_n326_));
  INV_X1    g125(.A(G148gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n324_), .A2(new_n328_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n331_), .B(new_n320_), .C1(new_n312_), .C2(new_n314_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n323_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(KEYINPUT29), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT78), .B(KEYINPUT28), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT79), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n334_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(G78gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G106gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n333_), .A2(KEYINPUT29), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n345_), .A2(new_n226_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G22gat), .B(G50gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n348_), .A3(new_n343_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  INV_X1    g154(.A(G134gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G127gat), .ZN(new_n357_));
  INV_X1    g156(.A(G127gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(G134gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n355_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n358_), .A2(G134gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n356_), .A2(G127gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT75), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n355_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n323_), .A2(new_n370_), .A3(new_n371_), .A4(new_n332_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n323_), .A2(new_n370_), .A3(new_n332_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT84), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT76), .A4(new_n368_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n363_), .A2(new_n369_), .A3(new_n376_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n375_), .A2(new_n377_), .B1(new_n323_), .B2(new_n332_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n354_), .B(new_n372_), .C1(new_n374_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n375_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT85), .B(KEYINPUT4), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n380_), .A2(new_n333_), .A3(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n372_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(KEYINPUT4), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n379_), .B1(new_n384_), .B2(new_n354_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G85gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT0), .B(G57gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n391_), .B(new_n379_), .C1(new_n384_), .C2(new_n354_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(KEYINPUT93), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT93), .B1(new_n390_), .B2(new_n392_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G15gat), .B(G43gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT74), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT30), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(new_n272_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G71gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n400_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n380_), .B(KEYINPUT31), .ZN(new_n404_));
  INV_X1    g203(.A(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n406_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n396_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n310_), .A2(new_n353_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT91), .B1(new_n305_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n390_), .A2(new_n392_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n282_), .A2(new_n283_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n413_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n418_));
  INV_X1    g217(.A(new_n413_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n299_), .B1(new_n301_), .B2(new_n295_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n420_), .A2(KEYINPUT90), .B1(new_n226_), .B2(new_n272_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n260_), .B1(new_n421_), .B2(new_n300_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n418_), .B(new_n419_), .C1(new_n422_), .C2(new_n292_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n384_), .A2(new_n354_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT88), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n384_), .A2(KEYINPUT88), .A3(new_n354_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n383_), .A2(KEYINPUT87), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n354_), .B1(new_n383_), .B2(KEYINPUT87), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n389_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n390_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n385_), .A2(new_n434_), .A3(new_n435_), .A4(new_n389_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n285_), .A2(new_n288_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n433_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n390_), .A2(new_n392_), .B1(new_n416_), .B2(new_n413_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(KEYINPUT92), .A3(new_n414_), .A4(new_n423_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n426_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n353_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n352_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n289_), .A2(new_n306_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n412_), .B1(new_n450_), .B2(new_n409_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n444_), .B2(new_n353_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n409_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n452_), .A2(KEYINPUT94), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n411_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n456_));
  INV_X1    g255(.A(G106gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n405_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n456_), .B(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT7), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G85gat), .B(G92gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT10), .B(G99gat), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n457_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n459_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(KEYINPUT65), .ZN(new_n474_));
  OR3_X1    g273(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT65), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT64), .B(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n474_), .B(new_n475_), .C1(new_n478_), .C2(KEYINPUT9), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G78gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT11), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(new_n482_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n483_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n468_), .A2(new_n480_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n468_), .B2(new_n480_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT12), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G230gat), .A2(G233gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n468_), .A2(new_n480_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n490_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n465_), .A2(new_n467_), .B1(new_n479_), .B2(new_n471_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n487_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n491_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G120gat), .B(G148gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT5), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G176gat), .B(G204gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n497_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n497_), .A2(KEYINPUT67), .A3(new_n502_), .A4(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n497_), .A2(new_n502_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n506_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n512_), .A2(KEYINPUT13), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT13), .B1(new_n512_), .B2(new_n514_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G29gat), .B(G36gat), .Z(new_n519_));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  INV_X1    g322(.A(G1gat), .ZN(new_n524_));
  INV_X1    g323(.A(G8gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G8gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n522_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n521_), .B(KEYINPUT15), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n529_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n529_), .B2(new_n522_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n533_), .B1(new_n536_), .B2(new_n532_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n537_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n518_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n455_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT36), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT69), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n498_), .A2(new_n521_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n552_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n492_), .A2(new_n534_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n558_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n551_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n492_), .A2(new_n522_), .B1(KEYINPUT35), .B2(new_n554_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n534_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n498_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n557_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n549_), .A2(KEYINPUT36), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n560_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n568_), .A2(KEYINPUT68), .A3(new_n560_), .A4(new_n569_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n546_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n529_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n493_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n580_), .B2(KEYINPUT17), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(KEYINPUT17), .B2(new_n577_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n580_), .A2(KEYINPUT70), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n550_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT37), .B1(new_n585_), .B2(new_n570_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n573_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n545_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n524_), .A3(new_n396_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n570_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n584_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n455_), .A2(new_n544_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n396_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n592_), .A2(new_n598_), .ZN(G1324gat));
  AOI21_X1  g398(.A(new_n525_), .B1(KEYINPUT97), .B2(KEYINPUT39), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n596_), .B2(new_n310_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n589_), .A2(new_n525_), .A3(new_n309_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(G1325gat));
  NOR4_X1   g407(.A1(new_n545_), .A2(G15gat), .A3(new_n409_), .A4(new_n588_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT99), .Z(new_n610_));
  INV_X1    g409(.A(new_n596_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n453_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n612_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(new_n612_), .B2(G15gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT100), .ZN(G1326gat));
  INV_X1    g415(.A(G22gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n589_), .A2(new_n617_), .A3(new_n352_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n611_), .B2(new_n352_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n624_), .B2(new_n625_), .ZN(G1327gat));
  INV_X1    g425(.A(new_n584_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n545_), .A2(new_n627_), .A3(new_n593_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n396_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n450_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT94), .B1(new_n452_), .B2(new_n453_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n309_), .A2(new_n352_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n630_), .A2(new_n631_), .B1(new_n632_), .B2(new_n410_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n573_), .A2(new_n586_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(new_n634_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n455_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n517_), .A2(new_n542_), .A3(new_n584_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT103), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n644_), .B(new_n641_), .C1(new_n635_), .C2(new_n638_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n396_), .A2(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n629_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  INV_X1    g447(.A(G36gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n628_), .A2(new_n649_), .A3(new_n309_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n643_), .A2(new_n645_), .A3(new_n310_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n653_), .B(KEYINPUT46), .C1(new_n654_), .C2(new_n649_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n654_), .A2(new_n649_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n652_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1329gat));
  AOI21_X1  g458(.A(G43gat), .B1(new_n628_), .B2(new_n453_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n453_), .A2(G43gat), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n646_), .B2(new_n665_), .ZN(new_n666_));
  NOR4_X1   g465(.A1(new_n643_), .A2(new_n645_), .A3(KEYINPUT105), .A4(new_n664_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT47), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n670_), .B(new_n662_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1330gat));
  NOR2_X1   g471(.A1(new_n353_), .A2(G50gat), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT108), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n628_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n646_), .A2(new_n352_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT107), .B1(new_n676_), .B2(G50gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(G1331gat));
  NAND2_X1  g478(.A1(new_n518_), .A2(new_n587_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT109), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n542_), .A3(new_n633_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n396_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n517_), .A2(new_n542_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n455_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n595_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT110), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n396_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n684_), .B1(new_n689_), .B2(new_n683_), .ZN(G1332gat));
  INV_X1    g489(.A(G64gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n691_), .A3(new_n309_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT48), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n309_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G64gat), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT48), .B(new_n691_), .C1(new_n688_), .C2(new_n309_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n682_), .A2(new_n698_), .A3(new_n453_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT49), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n688_), .A2(new_n453_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(G71gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT49), .B(new_n698_), .C1(new_n688_), .C2(new_n453_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1334gat));
  NAND3_X1  g503(.A1(new_n682_), .A2(new_n339_), .A3(new_n352_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n688_), .A2(new_n352_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G78gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT50), .B(new_n339_), .C1(new_n688_), .C2(new_n352_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1335gat));
  AND3_X1   g509(.A1(new_n686_), .A2(new_n584_), .A3(new_n594_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n396_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n685_), .A2(new_n584_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n597_), .A2(new_n476_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT111), .Z(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n714_), .B2(new_n716_), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n477_), .A3(new_n309_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n714_), .A2(new_n309_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n477_), .ZN(G1337gat));
  AOI21_X1  g519(.A(new_n405_), .B1(new_n714_), .B2(new_n453_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n453_), .A2(new_n469_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n711_), .B2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n711_), .A2(new_n457_), .A3(new_n352_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n714_), .A2(new_n352_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G106gat), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT52), .B(new_n457_), .C1(new_n714_), .C2(new_n352_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g531(.A(KEYINPUT118), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n512_), .A2(new_n542_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n497_), .B2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n489_), .A2(KEYINPUT12), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n500_), .B2(KEYINPUT12), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n491_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n495_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(new_n501_), .A3(new_n738_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n501_), .B1(new_n742_), .B2(new_n738_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(KEYINPUT55), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n506_), .B1(new_n741_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n490_), .A2(new_n496_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n736_), .B1(new_n749_), .B2(new_n501_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n737_), .B(new_n740_), .C1(new_n750_), .C2(new_n743_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n506_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n734_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n512_), .A2(new_n514_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n537_), .A2(new_n541_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n540_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT115), .Z(new_n757_));
  AOI21_X1  g556(.A(new_n531_), .B1(new_n536_), .B2(KEYINPUT116), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(KEYINPUT116), .B2(new_n536_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n754_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n593_), .B1(new_n753_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n734_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n506_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n506_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n761_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT57), .A3(new_n593_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n748_), .A2(new_n773_), .A3(new_n752_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n512_), .A2(new_n760_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n768_), .B2(KEYINPUT117), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n774_), .A2(KEYINPUT58), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT58), .B1(new_n774_), .B2(new_n776_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n634_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n584_), .B1(new_n772_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT13), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n754_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n512_), .A2(KEYINPUT13), .A3(new_n514_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n587_), .A2(new_n543_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT113), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n517_), .A2(new_n786_), .A3(new_n543_), .A4(new_n587_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(KEYINPUT54), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n784_), .A2(KEYINPUT113), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n597_), .B1(new_n780_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n632_), .A2(new_n453_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT59), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n767_), .A2(new_n768_), .A3(KEYINPUT117), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n746_), .A2(KEYINPUT117), .A3(new_n747_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n775_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n774_), .A2(new_n776_), .A3(KEYINPUT58), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n637_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n765_), .A3(new_n771_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n791_), .B1(new_n805_), .B2(new_n584_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  NOR4_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n597_), .A4(new_n794_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n733_), .B1(new_n796_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT57), .B1(new_n770_), .B2(new_n593_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n764_), .B(new_n594_), .C1(new_n769_), .C2(new_n761_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n627_), .B1(new_n812_), .B2(new_n804_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n396_), .B(new_n795_), .C1(new_n813_), .C2(new_n791_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n807_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n793_), .A2(KEYINPUT59), .A3(new_n795_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT118), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(new_n542_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G113gat), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n543_), .A2(G113gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n814_), .B2(new_n820_), .ZN(G1340gat));
  AOI21_X1  g620(.A(new_n517_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n822_));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n517_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(KEYINPUT60), .B2(new_n823_), .ZN(new_n825_));
  OAI22_X1  g624(.A1(new_n822_), .A2(new_n823_), .B1(new_n814_), .B2(new_n825_), .ZN(G1341gat));
  NOR2_X1   g625(.A1(new_n584_), .A2(new_n358_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n809_), .A2(new_n817_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n358_), .B1(new_n814_), .B2(new_n584_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(KEYINPUT119), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT119), .B1(new_n828_), .B2(new_n829_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1342gat));
  NAND4_X1  g631(.A1(new_n809_), .A2(G134gat), .A3(new_n817_), .A4(new_n637_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n814_), .A2(new_n593_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n834_), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT120), .B1(new_n834_), .B2(G134gat), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n833_), .A2(new_n835_), .A3(new_n836_), .ZN(G1343gat));
  NAND4_X1  g636(.A1(new_n793_), .A2(new_n352_), .A3(new_n409_), .A4(new_n310_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n543_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT121), .B(G141gat), .Z(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1344gat));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n517_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(new_n327_), .ZN(G1345gat));
  NOR2_X1   g642(.A1(new_n838_), .A2(new_n584_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT61), .B(G155gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  INV_X1    g645(.A(G162gat), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n838_), .A2(new_n847_), .A3(new_n634_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n838_), .B2(new_n593_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n850_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n806_), .A2(new_n310_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n396_), .A2(new_n352_), .A3(new_n409_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n543_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT123), .B(new_n854_), .C1(new_n858_), .C2(new_n234_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n234_), .B1(new_n860_), .B2(KEYINPUT62), .ZN(new_n861_));
  OAI221_X1 g660(.A(new_n861_), .B1(new_n860_), .B2(KEYINPUT62), .C1(new_n857_), .C2(new_n543_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT22), .B(G169gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n862_), .A3(new_n864_), .ZN(G1348gat));
  XOR2_X1   g664(.A(KEYINPUT124), .B(G176gat), .Z(new_n866_));
  NOR2_X1   g665(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n857_), .A2(new_n517_), .ZN(new_n868_));
  MUX2_X1   g667(.A(new_n866_), .B(new_n867_), .S(new_n868_), .Z(G1349gat));
  NAND4_X1  g668(.A1(new_n855_), .A2(new_n265_), .A3(new_n627_), .A4(new_n856_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT125), .Z(new_n871_));
  INV_X1    g670(.A(new_n857_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n627_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(G183gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(KEYINPUT126), .A3(new_n627_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n857_), .B2(new_n634_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n594_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n857_), .B2(new_n878_), .ZN(G1351gat));
  NOR3_X1   g678(.A1(new_n396_), .A2(new_n453_), .A3(new_n353_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n855_), .A2(new_n880_), .ZN(new_n881_));
  OAI22_X1  g680(.A1(new_n881_), .A2(new_n543_), .B1(KEYINPUT127), .B2(new_n212_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n212_), .A2(KEYINPUT127), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n882_), .B(new_n883_), .Z(G1352gat));
  NOR2_X1   g683(.A1(new_n881_), .A2(new_n517_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(G204gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n208_), .A2(new_n209_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1353gat));
  INV_X1    g687(.A(new_n881_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n627_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  AND2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n890_), .B2(new_n891_), .ZN(G1354gat));
  OR3_X1    g693(.A1(new_n881_), .A2(G218gat), .A3(new_n593_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G218gat), .B1(new_n881_), .B2(new_n634_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1355gat));
endmodule


