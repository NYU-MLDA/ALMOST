//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  OR3_X1    g000(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G183gat), .A3(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n209_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT76), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n202_), .A2(KEYINPUT24), .A3(new_n216_), .A4(new_n203_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n206_), .A2(new_n212_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n208_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT30), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G127gat), .B(G134gat), .Z(new_n229_));
  XOR2_X1   g028(.A(G113gat), .B(G120gat), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n231_), .A2(KEYINPUT79), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT79), .B1(new_n231_), .B2(new_n234_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n228_), .A2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(G15gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G71gat), .ZN(new_n244_));
  INV_X1    g043(.A(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT77), .B(G43gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT31), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n226_), .A2(new_n227_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n240_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n255_), .A2(new_n251_), .A3(new_n239_), .A4(new_n238_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G57gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT91), .Z(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT92), .Z(new_n264_));
  INV_X1    g063(.A(G141gat), .ZN(new_n265_));
  INV_X1    g064(.A(G148gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G155gat), .ZN(new_n276_));
  INV_X1    g075(.A(G162gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n275_), .A2(KEYINPUT1), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n279_), .A3(new_n274_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n270_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n268_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n276_), .A2(new_n277_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n288_), .A2(new_n275_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT81), .B1(new_n281_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n274_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT1), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n280_), .A3(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n269_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n288_), .A2(new_n275_), .A3(new_n289_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n299_), .A3(new_n237_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n281_), .A2(new_n290_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n231_), .A2(new_n234_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(new_n300_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n264_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n300_), .A2(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n263_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n261_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n310_), .A3(new_n261_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n257_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n316_));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n291_), .A2(new_n299_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n291_), .C2(new_n299_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n316_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n281_), .A2(new_n290_), .A3(KEYINPUT81), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n297_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n319_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT82), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n316_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G22gat), .B(G50gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n322_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT87), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n330_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n322_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT21), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G197gat), .ZN(new_n344_));
  INV_X1    g143(.A(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n340_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G211gat), .B(G218gat), .Z(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT85), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n350_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(KEYINPUT86), .A3(new_n340_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(new_n350_), .A3(new_n359_), .A4(KEYINPUT21), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n353_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n304_), .B2(new_n319_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(G228gat), .A3(G233gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n349_), .A2(new_n355_), .A3(new_n351_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(G228gat), .B2(G233gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n291_), .A2(KEYINPUT29), .A3(new_n299_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(KEYINPUT84), .B2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(KEYINPUT84), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G78gat), .B(G106gat), .Z(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n372_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n363_), .B(new_n374_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n333_), .A2(new_n339_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n336_), .A2(new_n338_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n378_), .A2(KEYINPUT87), .A3(new_n373_), .A4(new_n375_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  INV_X1    g180(.A(new_n208_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n219_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n209_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT89), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n212_), .B(new_n389_), .C1(G183gat), .C2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(G169gat), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n391_), .A2(KEYINPUT22), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(KEYINPUT22), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT88), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G169gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n388_), .A2(new_n390_), .A3(new_n400_), .A4(new_n216_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n205_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n217_), .A2(new_n215_), .A3(new_n220_), .A4(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n366_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n361_), .B2(new_n225_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT19), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n364_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n401_), .A2(new_n403_), .B1(new_n411_), .B2(new_n356_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n361_), .B2(new_n225_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n410_), .B1(new_n414_), .B2(new_n409_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G8gat), .B(G36gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT18), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n381_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n412_), .A2(new_n413_), .A3(new_n409_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n409_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n381_), .B(new_n420_), .C1(new_n422_), .C2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n404_), .A2(KEYINPUT90), .ZN(new_n426_));
  AOI211_X1 g225(.A(new_n405_), .B(new_n409_), .C1(new_n361_), .C2(new_n225_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n366_), .A2(new_n401_), .A3(new_n428_), .A4(new_n403_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n419_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT27), .B1(new_n421_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n420_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n432_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n315_), .A2(new_n380_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n314_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n257_), .B1(new_n380_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n430_), .A2(new_n443_), .A3(new_n431_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n264_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n300_), .A2(new_n306_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT4), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n450_), .B2(new_n302_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n309_), .A2(new_n263_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n261_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n447_), .B1(new_n454_), .B2(new_n311_), .ZN(new_n455_));
  OR2_X1    g254(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n308_), .A2(new_n310_), .A3(new_n261_), .A4(new_n456_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n263_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n261_), .B1(new_n309_), .B2(new_n264_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n458_), .A2(new_n436_), .A3(new_n432_), .A4(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n455_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n379_), .B2(new_n377_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n440_), .B1(new_n442_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT71), .ZN(new_n469_));
  INV_X1    g268(.A(G36gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G29gat), .ZN(new_n471_));
  INV_X1    g270(.A(G29gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G36gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT71), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT72), .B1(new_n469_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n473_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n468_), .A2(KEYINPUT71), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n475_), .A2(new_n483_), .A3(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  INV_X1    g287(.A(G1gat), .ZN(new_n489_));
  INV_X1    g288(.A(G8gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  NAND2_X1  g293(.A1(new_n487_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n487_), .A2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n467_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499_));
  INV_X1    g298(.A(new_n486_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n483_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n485_), .A2(KEYINPUT15), .A3(new_n486_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n495_), .B1(new_n504_), .B2(new_n494_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n505_), .B2(new_n467_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n506_), .B(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n465_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n245_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT65), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n516_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(KEYINPUT65), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT6), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(G99gat), .A3(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n524_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G85gat), .B(G92gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT8), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n530_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(KEYINPUT67), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n527_), .A2(new_n529_), .A3(KEYINPUT68), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n524_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n533_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n532_), .A2(new_n537_), .B1(new_n543_), .B2(KEYINPUT8), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(KEYINPUT9), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(G85gat), .A3(G92gat), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n530_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT10), .B(G99gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT64), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n515_), .B2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n544_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n514_), .B1(new_n504_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT34), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n552_), .A2(new_n487_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n502_), .B(new_n503_), .C1(new_n544_), .C2(new_n551_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT74), .ZN(new_n563_));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n558_), .A2(new_n561_), .B1(KEYINPUT36), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n556_), .B1(new_n560_), .B2(new_n514_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n560_), .B(new_n559_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n567_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n513_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n568_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT37), .A3(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n550_), .A2(new_n515_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(new_n530_), .A3(new_n545_), .A4(new_n547_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT11), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(KEYINPUT11), .ZN(new_n586_));
  XOR2_X1   g385(.A(G71gat), .B(G78gat), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n521_), .A2(new_n523_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n534_), .B1(new_n591_), .B2(new_n525_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n531_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT8), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n583_), .B(new_n590_), .C1(new_n593_), .C2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT12), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n543_), .A2(KEYINPUT8), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n531_), .B2(new_n592_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n590_), .B1(new_n599_), .B2(new_n583_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  INV_X1    g401(.A(new_n590_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n602_), .B(new_n603_), .C1(new_n544_), .C2(new_n551_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n581_), .B1(new_n601_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n544_), .B2(new_n551_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT69), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n596_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n581_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n609_), .B(new_n610_), .C1(new_n608_), .C2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n606_), .A2(new_n611_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT13), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n494_), .B(new_n590_), .Z(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626_));
  XOR2_X1   g425(.A(G127gat), .B(G155gat), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT16), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n625_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(KEYINPUT17), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n580_), .A2(new_n622_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n512_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT95), .ZN(new_n638_));
  INV_X1    g437(.A(new_n314_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n638_), .A2(G1gat), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT98), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n577_), .A2(new_n578_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT97), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n465_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n511_), .A3(new_n634_), .A4(new_n622_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n639_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n643_), .B(new_n648_), .C1(new_n641_), .C2(new_n640_), .ZN(G1324gat));
  OAI21_X1  g448(.A(G8gat), .B1(new_n647_), .B2(new_n439_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT39), .ZN(new_n651_));
  INV_X1    g450(.A(new_n439_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n490_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n638_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n647_), .B2(new_n257_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n257_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n242_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n658_), .B(new_n659_), .C1(new_n637_), .C2(new_n661_), .ZN(G1326gat));
  OAI21_X1  g461(.A(G22gat), .B1(new_n647_), .B2(new_n380_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT42), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n380_), .A2(G22gat), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT100), .Z(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n637_), .B2(new_n666_), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n644_), .A2(new_n634_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n512_), .A2(new_n622_), .A3(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT105), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n314_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n575_), .A2(new_n579_), .A3(KEYINPUT102), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT102), .B1(new_n575_), .B2(new_n579_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n465_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT43), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n580_), .A2(KEYINPUT43), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n465_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n465_), .A2(new_n677_), .A3(KEYINPUT103), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n634_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n622_), .A2(new_n511_), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT101), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(KEYINPUT44), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n686_), .B(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n639_), .A2(new_n472_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n671_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  NAND3_X1  g491(.A1(new_n670_), .A2(new_n470_), .A3(new_n652_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT45), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n689_), .A2(new_n439_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n470_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n694_), .B(new_n698_), .C1(new_n470_), .C2(new_n695_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  NOR2_X1   g501(.A1(new_n257_), .A2(G43gat), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n670_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n690_), .A2(new_n660_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G43gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n689_), .B2(new_n380_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n380_), .A2(G50gat), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT107), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n670_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n622_), .A2(new_n511_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n465_), .A2(new_n713_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(new_n634_), .A3(new_n580_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n314_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n646_), .A2(new_n634_), .A3(new_n713_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n639_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n718_), .B2(new_n439_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n439_), .A2(G64gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT109), .Z(new_n725_));
  NAND2_X1  g524(.A1(new_n715_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n718_), .B2(new_n257_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n715_), .A2(new_n731_), .A3(new_n660_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n718_), .B2(new_n380_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  INV_X1    g535(.A(new_n380_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n715_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1335gat));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n676_), .A2(new_n680_), .A3(new_n741_), .A4(new_n681_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n622_), .A2(new_n511_), .A3(new_n634_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT113), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(KEYINPUT43), .A2(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n741_), .B1(new_n746_), .B2(new_n681_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n740_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n682_), .A2(KEYINPUT112), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n749_), .A2(KEYINPUT114), .A3(new_n744_), .A4(new_n742_), .ZN(new_n750_));
  AND4_X1   g549(.A1(G85gat), .A2(new_n748_), .A3(new_n314_), .A4(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n714_), .A2(new_n668_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n314_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT111), .Z(new_n754_));
  OR2_X1    g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT115), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n752_), .B2(new_n652_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n748_), .A2(new_n750_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n652_), .A2(G92gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT116), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n759_), .B2(new_n761_), .ZN(G1337gat));
  NAND3_X1  g561(.A1(new_n752_), .A2(new_n660_), .A3(new_n550_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n748_), .A2(new_n660_), .A3(new_n750_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n764_), .A2(KEYINPUT117), .A3(G99gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT117), .B1(new_n764_), .B2(G99gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT51), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n763_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1338gat));
  AND2_X1   g570(.A1(new_n744_), .A2(new_n737_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n515_), .B1(new_n772_), .B2(new_n682_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT52), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n752_), .A2(new_n515_), .A3(new_n737_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g576(.A(new_n511_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n636_), .A2(KEYINPUT118), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n635_), .B2(new_n511_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(KEYINPUT54), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n780_), .B(new_n783_), .C1(new_n635_), .C2(new_n511_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n607_), .A2(KEYINPUT12), .A3(new_n596_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n610_), .A3(new_n604_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n610_), .B1(new_n787_), .B2(new_n604_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n581_), .C1(new_n601_), .C2(new_n605_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT120), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n606_), .A2(KEYINPUT55), .A3(new_n788_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT120), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n793_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n619_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n786_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n796_), .A2(new_n797_), .A3(new_n793_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n797_), .B1(new_n796_), .B2(new_n793_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n617_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n511_), .A2(KEYINPUT119), .A3(new_n620_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT119), .B1(new_n511_), .B2(new_n620_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n801_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n506_), .A2(new_n510_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n496_), .A2(new_n497_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n509_), .B1(new_n811_), .B2(new_n466_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n466_), .B1(new_n505_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n813_), .B2(new_n505_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n810_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n621_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n809_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT57), .A3(new_n644_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT123), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n644_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n644_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT57), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n816_), .A2(new_n620_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n804_), .B2(KEYINPUT56), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n799_), .A2(new_n786_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n580_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n804_), .A2(KEYINPUT56), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n799_), .A2(new_n786_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(KEYINPUT58), .A4(new_n829_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n833_), .A3(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n820_), .A2(new_n823_), .A3(new_n827_), .A4(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n785_), .B1(new_n838_), .B2(new_n683_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n737_), .A2(new_n652_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n314_), .A3(new_n660_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n511_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n841_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n837_), .B1(new_n825_), .B2(KEYINPUT57), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n826_), .B1(new_n825_), .B2(KEYINPUT57), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n634_), .B1(new_n850_), .B2(new_n827_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT59), .B(new_n847_), .C1(new_n851_), .C2(new_n785_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n778_), .B1(new_n846_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n844_), .B1(new_n853_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n842_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n622_), .B1(new_n846_), .B2(new_n852_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n842_), .A2(new_n860_), .A3(new_n634_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n683_), .B1(new_n846_), .B2(new_n852_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n846_), .A2(new_n852_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n833_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n842_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n645_), .A2(G134gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT124), .B1(new_n866_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n580_), .B1(new_n846_), .B2(new_n852_), .ZN(new_n872_));
  OAI221_X1 g671(.A(new_n871_), .B1(new_n867_), .B2(new_n868_), .C1(new_n872_), .C2(new_n864_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n380_), .A2(new_n660_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n876_), .A2(new_n639_), .A3(new_n652_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n839_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n511_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NOR3_X1   g680(.A1(new_n839_), .A2(new_n622_), .A3(new_n878_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT125), .B(G148gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n634_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT126), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n879_), .A2(new_n887_), .A3(new_n634_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1346gat));
  OR3_X1    g691(.A1(new_n839_), .A2(new_n645_), .A3(new_n878_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n672_), .A2(new_n673_), .A3(new_n277_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n893_), .A2(new_n277_), .B1(new_n879_), .B2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n839_), .A2(new_n439_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n315_), .A2(new_n380_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n511_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n896_), .A2(new_n511_), .A3(new_n398_), .A4(new_n897_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1348gat));
  NAND2_X1  g702(.A1(new_n896_), .A2(new_n897_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n622_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n399_), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n896_), .A2(new_n634_), .A3(new_n897_), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n213_), .B(G183gat), .S(new_n907_), .Z(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n904_), .B2(new_n580_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n214_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n645_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n904_), .B2(new_n911_), .ZN(G1351gat));
  NOR2_X1   g711(.A1(new_n876_), .A2(new_n314_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n896_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n778_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n344_), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n914_), .A2(new_n622_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n345_), .ZN(G1353gat));
  AOI21_X1  g717(.A(new_n683_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n896_), .A2(new_n913_), .A3(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n920_), .B(new_n922_), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n914_), .B2(new_n580_), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n645_), .A2(G218gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n914_), .B2(new_n925_), .ZN(G1355gat));
endmodule


