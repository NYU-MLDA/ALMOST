//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202_));
  XOR2_X1   g001(.A(G190gat), .B(G218gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G85gat), .B(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n207_), .A2(G85gat), .A3(G92gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT8), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n206_), .B1(new_n219_), .B2(KEYINPUT8), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n218_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n218_), .B2(new_n222_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n215_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G29gat), .B(G36gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G43gat), .B(G50gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n227_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT15), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n218_), .A2(new_n222_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n221_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n218_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n231_), .A3(new_n215_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT34), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n239_), .A2(new_n215_), .B1(new_n232_), .B2(new_n230_), .ZN(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT35), .B(new_n243_), .C1(new_n244_), .C2(KEYINPUT68), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n243_), .A2(KEYINPUT35), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n241_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n225_), .B2(new_n233_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT35), .ZN(new_n250_));
  INV_X1    g049(.A(new_n243_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n241_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n202_), .B(new_n205_), .C1(new_n248_), .C2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n252_), .B2(new_n246_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n205_), .A2(new_n202_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n205_), .A2(new_n202_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n245_), .A2(new_n241_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT22), .B(G169gat), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT82), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n269_));
  OAI211_X1 g068(.A(KEYINPUT82), .B(new_n266_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n264_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n281_), .B2(KEYINPUT23), .ZN(new_n282_));
  INV_X1    g081(.A(G183gat), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n283_), .A2(KEYINPUT79), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(KEYINPUT79), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT80), .B(G190gat), .Z(new_n287_));
  OAI21_X1  g086(.A(new_n282_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT83), .B(new_n264_), .C1(new_n267_), .C2(new_n271_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n274_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(KEYINPUT25), .A3(new_n285_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT25), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G190gat), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n294_), .B(new_n296_), .C1(new_n295_), .C2(new_n287_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT24), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n297_), .A2(new_n300_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n290_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT30), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G71gat), .B(G99gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(KEYINPUT30), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G43gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n313_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n306_), .B(KEYINPUT30), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n308_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n318_), .B2(new_n311_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n263_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n313_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n316_), .A3(new_n311_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n321_), .A2(G227gat), .A3(G233gat), .A4(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n323_), .A3(KEYINPUT84), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT31), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n320_), .A2(new_n323_), .A3(KEYINPUT84), .A4(new_n328_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT89), .B(G197gat), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT21), .B(new_n334_), .C1(new_n335_), .C2(G204gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G197gat), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n339_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT90), .B1(new_n339_), .B2(G204gat), .ZN(new_n341_));
  INV_X1    g140(.A(G204gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n340_), .B(new_n341_), .C1(new_n335_), .C2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n336_), .B(new_n338_), .C1(new_n343_), .C2(KEYINPUT21), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(KEYINPUT21), .A3(new_n337_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT86), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(new_n347_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT2), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n347_), .B1(new_n358_), .B2(KEYINPUT1), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n355_), .A3(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n346_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT88), .Z(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n346_), .B2(KEYINPUT91), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G78gat), .B(G106gat), .Z(new_n373_));
  OAI221_X1 g172(.A(new_n346_), .B1(KEYINPUT91), .B2(new_n370_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n333_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n376_), .A2(new_n333_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n366_), .A2(new_n367_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n379_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n377_), .A2(new_n378_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT92), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT92), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n388_), .B(new_n383_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  INV_X1    g193(.A(new_n282_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT94), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n293_), .A2(new_n400_), .A3(new_n396_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G190gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT26), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n296_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n304_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n395_), .B1(new_n408_), .B2(KEYINPUT95), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n304_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n302_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n283_), .A2(new_n403_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n298_), .A2(new_n299_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n416_), .A2(new_n417_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n298_), .A2(KEYINPUT96), .A3(new_n299_), .A4(new_n415_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(new_n264_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n409_), .A2(new_n414_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n344_), .A2(new_n345_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n394_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI211_X1 g222(.A(KEYINPUT97), .B(new_n422_), .C1(new_n290_), .C2(new_n305_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n306_), .B2(new_n346_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n393_), .B(new_n423_), .C1(new_n424_), .C2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G92gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT18), .B(G64gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT32), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n421_), .A2(new_n422_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n290_), .A2(new_n305_), .A3(new_n422_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT20), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n392_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n327_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n361_), .A2(new_n365_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(KEYINPUT99), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT99), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n361_), .A2(new_n441_), .A3(new_n365_), .A4(new_n327_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(KEYINPUT4), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n439_), .A2(KEYINPUT100), .A3(new_n446_), .A4(new_n438_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n439_), .A2(new_n446_), .A3(new_n438_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT100), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .A4(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n440_), .A2(new_n442_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n444_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT0), .B(G57gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n451_), .A2(new_n453_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n437_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n423_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n392_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n435_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n393_), .C1(new_n422_), .C2(new_n421_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n432_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT102), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n412_), .A2(new_n413_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT95), .B1(new_n410_), .B2(new_n411_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n282_), .A3(new_n303_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n420_), .A2(new_n418_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n422_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT20), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n306_), .A2(new_n346_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT97), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n306_), .A2(new_n425_), .A3(new_n346_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n466_), .B1(new_n478_), .B2(new_n393_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n432_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n451_), .A2(new_n453_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n458_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n451_), .A2(new_n453_), .A3(new_n459_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT102), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n481_), .A2(new_n485_), .A3(new_n486_), .A4(new_n437_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n468_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n443_), .A2(new_n444_), .A3(new_n447_), .A4(new_n450_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n452_), .B(KEYINPUT101), .Z(new_n490_));
  OAI211_X1 g289(.A(new_n458_), .B(new_n489_), .C1(new_n490_), .C2(new_n444_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n484_), .B(KEYINPUT33), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n427_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n431_), .B1(new_n427_), .B2(new_n436_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT98), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n427_), .A2(new_n436_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT98), .ZN(new_n497_));
  INV_X1    g296(.A(new_n431_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n491_), .B(new_n492_), .C1(new_n495_), .C2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n390_), .B1(new_n488_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n485_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n498_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n427_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n497_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n493_), .B1(new_n494_), .B2(KEYINPUT98), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n479_), .A2(new_n498_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT27), .A3(new_n504_), .ZN(new_n510_));
  AND4_X1   g309(.A1(new_n502_), .A2(new_n508_), .A3(new_n390_), .A4(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n332_), .B1(new_n501_), .B2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n508_), .A2(new_n513_), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT103), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n330_), .A2(new_n331_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT103), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n508_), .A2(new_n513_), .A3(new_n517_), .A4(new_n510_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n502_), .A4(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n262_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n225_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n215_), .B(new_n529_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT12), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n225_), .A2(new_n534_), .A3(new_n530_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n522_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n521_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G176gat), .B(G204gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G120gat), .B(G148gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  NOR3_X1   g341(.A1(new_n536_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(KEYINPUT13), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(KEYINPUT13), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G15gat), .B(G22gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT70), .B(G1gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G8gat), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n555_), .B2(KEYINPUT14), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G1gat), .B(G8gat), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n231_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n557_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n555_), .A2(KEYINPUT14), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n553_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n557_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n228_), .A3(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n560_), .A2(KEYINPUT74), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT74), .B1(new_n560_), .B2(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n552_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT75), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n558_), .A2(new_n559_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n233_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT76), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n233_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n551_), .A3(new_n560_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n558_), .A2(new_n559_), .A3(new_n231_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n228_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n560_), .A2(KEYINPUT74), .A3(new_n565_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n552_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n569_), .A2(new_n575_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n339_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT77), .B(G169gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n569_), .A2(new_n575_), .A3(new_n583_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n550_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT72), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n529_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n570_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n603_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n593_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n520_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n502_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT78), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n592_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT69), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n255_), .A2(new_n260_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n255_), .B2(new_n260_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n261_), .A2(KEYINPUT69), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n255_), .A2(new_n260_), .A3(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT37), .A3(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n607_), .B(KEYINPUT73), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n550_), .B(KEYINPUT67), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n616_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n485_), .B(KEYINPUT104), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n630_), .A2(new_n554_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n612_), .B1(new_n638_), .B2(new_n639_), .ZN(G1324gat));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n512_), .A2(new_n519_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n508_), .A2(new_n510_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n261_), .A4(new_n609_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT106), .B1(new_n644_), .B2(G8gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n644_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(KEYINPUT107), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n652_), .A3(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(new_n643_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n630_), .A2(G8gat), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n641_), .B(new_n656_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n653_), .A2(KEYINPUT40), .A3(new_n655_), .A4(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n611_), .B2(new_n332_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n630_), .A2(G15gat), .A3(new_n332_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n610_), .B2(new_n390_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT42), .Z(new_n669_));
  NAND2_X1  g468(.A1(new_n390_), .A2(new_n667_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n630_), .B2(new_n670_), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n621_), .A2(new_n624_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(KEYINPUT43), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n642_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n621_), .A2(new_n624_), .A3(KEYINPUT109), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n680_));
  OAI21_X1  g479(.A(new_n674_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n593_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n626_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n682_), .A4(new_n626_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n685_), .A2(G29gat), .A3(new_n631_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G29gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n626_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n261_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n616_), .A2(new_n550_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n691_), .B2(new_n502_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n687_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT110), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n695_), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n686_), .A2(new_n643_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n685_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n691_), .A2(G36gat), .A3(new_n654_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n702_), .A2(KEYINPUT45), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(KEYINPUT45), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n683_), .A2(new_n684_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n686_), .A2(new_n643_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G36gat), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(KEYINPUT46), .A3(new_n703_), .A4(new_n704_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n691_), .B2(new_n332_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n686_), .A2(G43gat), .A3(new_n516_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n707_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g515(.A1(new_n686_), .A2(new_n390_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G50gat), .B1(new_n707_), .B2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n513_), .A2(G50gat), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT111), .Z(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n691_), .B2(new_n720_), .ZN(G1331gat));
  NOR2_X1   g520(.A1(new_n614_), .A2(new_n626_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n520_), .A2(new_n628_), .A3(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT112), .B(G57gat), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n723_), .A2(new_n502_), .A3(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n550_), .A2(new_n592_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n642_), .A2(new_n627_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n631_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1332gat));
  OAI21_X1  g528(.A(G64gat), .B1(new_n723_), .B2(new_n654_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT48), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n654_), .A2(G64gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT113), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n727_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n727_), .A2(new_n736_), .A3(new_n516_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n738_));
  INV_X1    g537(.A(new_n723_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n516_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(G71gat), .ZN(new_n741_));
  AOI211_X1 g540(.A(KEYINPUT49), .B(new_n736_), .C1(new_n739_), .C2(new_n516_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n737_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT114), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n723_), .B2(new_n513_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n727_), .A2(new_n747_), .A3(new_n390_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1335gat));
  INV_X1    g548(.A(new_n592_), .ZN(new_n750_));
  AND4_X1   g549(.A1(new_n642_), .A2(new_n750_), .A3(new_n628_), .A4(new_n690_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n631_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n726_), .A2(new_n626_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n681_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n502_), .A2(new_n455_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n751_), .B2(new_n643_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n643_), .A2(G92gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n755_), .B2(new_n759_), .ZN(G1337gat));
  NAND3_X1  g559(.A1(new_n681_), .A2(new_n516_), .A3(new_n754_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G99gat), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n516_), .A2(new_n209_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n751_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n762_), .A2(new_n764_), .B1(KEYINPUT115), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(KEYINPUT115), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n681_), .A2(new_n390_), .A3(new_n754_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G106gat), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n751_), .A2(new_n210_), .A3(new_n390_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n771_), .A2(new_n772_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n769_), .A2(G106gat), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n774_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n773_), .A2(new_n780_), .A3(new_n774_), .A4(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n722_), .A2(new_n550_), .A3(new_n672_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n783_), .B(new_n784_), .Z(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n533_), .A2(new_n522_), .A3(new_n535_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n533_), .A2(new_n535_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n521_), .ZN(new_n790_));
  AOI211_X1 g589(.A(KEYINPUT55), .B(new_n522_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n542_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n581_), .A2(new_n551_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n572_), .A2(new_n552_), .A3(new_n560_), .A4(new_n574_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n588_), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n591_), .A2(KEYINPUT120), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT120), .B1(new_n591_), .B2(new_n797_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n794_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n792_), .A2(new_n802_), .A3(new_n542_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n544_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n786_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n804_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n800_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n798_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n806_), .A2(new_n808_), .A3(KEYINPUT58), .A4(new_n794_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n625_), .A2(new_n805_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n547_), .B1(new_n807_), .B2(new_n798_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n592_), .B2(new_n544_), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT118), .B(new_n543_), .C1(new_n589_), .C2(new_n591_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n802_), .A2(KEYINPUT119), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n792_), .A2(new_n542_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n792_), .B2(new_n542_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n811_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT57), .B1(new_n820_), .B2(new_n262_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n592_), .A2(new_n544_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT118), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n592_), .A2(new_n812_), .A3(new_n544_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n819_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n811_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n261_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n810_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n785_), .B1(new_n607_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n632_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n592_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n830_), .B2(new_n689_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n625_), .A2(new_n805_), .A3(new_n809_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n828_), .B1(new_n827_), .B2(new_n261_), .ZN(new_n840_));
  AOI211_X1 g639(.A(KEYINPUT57), .B(new_n262_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(KEYINPUT121), .A3(new_n626_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n838_), .A2(new_n843_), .A3(new_n785_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n833_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n783_), .B(new_n784_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n608_), .B2(new_n842_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n833_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n614_), .A2(G113gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n836_), .B1(new_n851_), .B2(new_n852_), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n628_), .A3(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT123), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n846_), .A2(new_n856_), .A3(new_n628_), .A4(new_n850_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(G120gat), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n550_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(G120gat), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT122), .B1(new_n860_), .B2(G120gat), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n835_), .B(new_n863_), .C1(new_n861_), .C2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n858_), .A2(new_n865_), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n834_), .B2(new_n626_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AND4_X1   g669(.A1(G127gat), .A2(new_n846_), .A3(new_n607_), .A4(new_n850_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n868_), .A2(new_n869_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(G1342gat));
  AOI21_X1  g672(.A(G134gat), .B1(new_n835_), .B2(new_n262_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n625_), .A2(G134gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n851_), .B2(new_n875_), .ZN(G1343gat));
  NAND4_X1  g675(.A1(new_n332_), .A2(new_n390_), .A3(new_n654_), .A4(new_n631_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT125), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n848_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n592_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT126), .B(G141gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n628_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n689_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  AOI21_X1  g686(.A(G162gat), .B1(new_n879_), .B2(new_n262_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n676_), .A2(G162gat), .A3(new_n677_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n879_), .B2(new_n889_), .ZN(G1347gat));
  NOR3_X1   g689(.A1(new_n332_), .A2(new_n654_), .A3(new_n631_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n844_), .A2(new_n513_), .A3(new_n592_), .A4(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G169gat), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n265_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n894_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n893_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1348gat));
  NAND3_X1  g699(.A1(new_n844_), .A2(new_n513_), .A3(new_n891_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902_), .B2(new_n859_), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n848_), .A2(new_n266_), .A3(new_n390_), .A4(new_n629_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n891_), .B2(new_n904_), .ZN(G1349gat));
  NOR3_X1   g704(.A1(new_n901_), .A2(new_n402_), .A3(new_n608_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n286_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n831_), .A2(new_n513_), .A3(new_n689_), .A4(new_n891_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n901_), .B2(new_n672_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n262_), .A2(new_n406_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n901_), .B2(new_n911_), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n654_), .A2(new_n485_), .A3(new_n513_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n831_), .A2(new_n332_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n831_), .A2(KEYINPUT127), .A3(new_n332_), .A4(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n592_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G197gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n918_), .A2(new_n339_), .A3(new_n592_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1352gat));
  AOI21_X1  g721(.A(G204gat), .B1(new_n918_), .B2(new_n628_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n342_), .B(new_n629_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  OR2_X1    g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n918_), .B2(new_n607_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT63), .B(G211gat), .ZN(new_n928_));
  AOI211_X1 g727(.A(new_n608_), .B(new_n928_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1354gat));
  AOI21_X1  g729(.A(G218gat), .B1(new_n918_), .B2(new_n262_), .ZN(new_n931_));
  INV_X1    g730(.A(G218gat), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n932_), .B(new_n672_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1355gat));
endmodule


