//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT75), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n206_), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n203_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT76), .ZN(new_n210_));
  XOR2_X1   g009(.A(G1gat), .B(G8gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n212_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G229gat), .A2(G233gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n222_), .B(new_n218_), .C1(new_n216_), .C2(new_n212_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT77), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n228_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G85gat), .B(G92gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT68), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT6), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT7), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(KEYINPUT66), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n239_), .ZN(new_n243_));
  OAI221_X1 g042(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .C1(new_n243_), .C2(KEYINPUT67), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n235_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n247_));
  NAND2_X1  g046(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n248_), .B(new_n235_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT10), .B(G99gat), .Z(new_n251_));
  INV_X1    g050(.A(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT9), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(G85gat), .A3(G92gat), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n237_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n234_), .A2(KEYINPUT9), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(KEYINPUT65), .A3(new_n252_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n250_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G57gat), .B(G64gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT11), .ZN(new_n266_));
  XOR2_X1   g065(.A(G71gat), .B(G78gat), .Z(new_n267_));
  OR2_X1    g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n263_), .B(KEYINPUT70), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n271_), .A3(new_n267_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n262_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n261_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n278_));
  OAI22_X1  g077(.A1(new_n278_), .A2(new_n273_), .B1(KEYINPUT72), .B2(KEYINPUT12), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G230gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT64), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n278_), .A2(new_n273_), .B1(KEYINPUT72), .B2(KEYINPUT12), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n282_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n262_), .B2(new_n274_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n278_), .B2(new_n273_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n262_), .A2(new_n288_), .A3(new_n274_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n287_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n280_), .A2(KEYINPUT73), .A3(new_n282_), .A4(new_n283_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n286_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G120gat), .B(G148gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT5), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G176gat), .B(G204gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n286_), .A2(new_n292_), .A3(new_n293_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT13), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(KEYINPUT13), .A3(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT31), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n309_), .A2(new_n310_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n310_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n312_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n313_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G169gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT23), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(G183gat), .A3(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n323_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n327_), .A2(KEYINPUT81), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n326_), .B2(KEYINPUT23), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n329_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  OR3_X1    g135(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT26), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G190gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT78), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n349_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n348_), .B1(new_n354_), .B2(KEYINPUT79), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n350_), .A2(KEYINPUT78), .ZN(new_n357_));
  OAI21_X1  g156(.A(G183gat), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n349_), .A2(KEYINPUT25), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT79), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n343_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n338_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI211_X1 g163(.A(KEYINPUT80), .B(new_n343_), .C1(new_n355_), .C2(new_n361_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n332_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  INV_X1    g166(.A(G43gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G227gat), .A2(G233gat), .ZN(new_n371_));
  INV_X1    g170(.A(G15gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT30), .ZN(new_n374_));
  INV_X1    g173(.A(new_n369_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n332_), .B(new_n375_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n370_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n374_), .B1(new_n370_), .B2(new_n376_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT84), .B(new_n320_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n336_), .A2(new_n337_), .ZN(new_n381_));
  OAI211_X1 g180(.A(KEYINPUT79), .B(G183gat), .C1(new_n356_), .C2(new_n357_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT26), .B(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n359_), .A2(KEYINPUT79), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n354_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n342_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n387_), .B2(KEYINPUT80), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n362_), .A2(new_n363_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n375_), .B1(new_n390_), .B2(new_n332_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n376_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n380_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n370_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n312_), .A4(new_n317_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n394_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT84), .B1(new_n397_), .B2(new_n320_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  AND2_X1   g207(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n409_));
  NOR2_X1   g208(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT2), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT2), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n417_));
  INV_X1    g216(.A(G141gat), .ZN(new_n418_));
  INV_X1    g217(.A(G148gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n416_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n413_), .A2(new_n415_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT87), .A3(new_n411_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n407_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(new_n412_), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n406_), .B(KEYINPUT1), .Z(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(new_n405_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT88), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n407_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT87), .B1(new_n425_), .B2(new_n411_), .ZN(new_n433_));
  AND4_X1   g232(.A1(KEYINPUT87), .A2(new_n411_), .A3(new_n416_), .A4(new_n421_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n436_));
  INV_X1    g235(.A(new_n430_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n402_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n402_), .A3(new_n440_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n401_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI211_X1 g243(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n431_), .C2(new_n438_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n441_), .A2(new_n445_), .A3(new_n400_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT21), .ZN(new_n447_));
  INV_X1    g246(.A(G204gat), .ZN(new_n448_));
  INV_X1    g247(.A(G197gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT89), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G197gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G197gat), .A2(G204gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n447_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G218gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G211gat), .ZN(new_n457_));
  INV_X1    g256(.A(G211gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G218gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(new_n452_), .A3(new_n448_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n447_), .B1(G197gat), .B2(G204gat), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n453_), .A2(new_n454_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT21), .A3(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(G228gat), .B2(G233gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G78gat), .B(G106gat), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n464_), .A2(new_n466_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n440_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n477_));
  OAI211_X1 g276(.A(G228gat), .B(G233gat), .C1(new_n476_), .C2(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n470_), .A2(new_n472_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n472_), .B1(new_n470_), .B2(new_n478_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n444_), .A2(new_n446_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n442_), .A2(new_n443_), .A3(new_n401_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n400_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n470_), .A2(new_n472_), .A3(new_n478_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n399_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G225gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n309_), .B(KEYINPUT82), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n431_), .A2(new_n438_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n435_), .A2(new_n309_), .A3(new_n437_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT4), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n494_), .B1(new_n499_), .B2(new_n490_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G1gat), .B(G29gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G85gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT0), .B(G57gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n492_), .A2(new_n493_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT4), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n490_), .A3(new_n496_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n494_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n504_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT27), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G226gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(new_n467_), .B(new_n331_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n323_), .B1(new_n336_), .B2(new_n325_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT25), .B(G183gat), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n383_), .A2(new_n521_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n330_), .A2(KEYINPUT92), .A3(new_n337_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT92), .B1(new_n330_), .B2(new_n337_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n527_), .A2(KEYINPUT93), .A3(new_n523_), .A4(new_n522_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n519_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT20), .B1(new_n529_), .B2(new_n468_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n517_), .B1(new_n518_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G8gat), .B(G36gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT18), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G64gat), .B(G92gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n366_), .A2(new_n467_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n468_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT20), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n517_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n531_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n535_), .B1(new_n531_), .B2(new_n540_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n514_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n535_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n518_), .A2(new_n530_), .A3(new_n517_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n517_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n524_), .A2(new_n525_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(new_n519_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n476_), .B2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n546_), .B1(new_n549_), .B2(new_n536_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n544_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n531_), .A2(new_n540_), .A3(new_n535_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT27), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT96), .B1(new_n543_), .B2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n543_), .A2(new_n553_), .A3(KEYINPUT96), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n488_), .B(new_n513_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT97), .ZN(new_n557_));
  INV_X1    g356(.A(new_n554_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n543_), .A2(new_n553_), .A3(KEYINPUT96), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n513_), .A4(new_n488_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n497_), .A2(new_n498_), .A3(new_n489_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT33), .B(new_n511_), .C1(new_n564_), .C2(new_n494_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n526_), .A2(new_n528_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n519_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n538_), .B1(new_n570_), .B2(new_n467_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n390_), .A2(new_n468_), .A3(new_n332_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n546_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n537_), .A2(new_n539_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n468_), .B1(new_n390_), .B2(new_n332_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n544_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n552_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n504_), .B1(new_n506_), .B2(new_n489_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n507_), .A2(new_n496_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n489_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n510_), .A2(KEYINPUT94), .A3(KEYINPUT33), .A4(new_n511_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n567_), .A2(new_n582_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(KEYINPUT32), .B(new_n535_), .C1(new_n545_), .C2(new_n550_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n535_), .A2(KEYINPUT32), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n531_), .A2(new_n540_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n587_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n589_), .B(new_n592_), .C1(new_n505_), .C2(new_n512_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n487_), .B1(new_n586_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n513_), .A2(new_n487_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n543_), .A2(new_n553_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n399_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n233_), .B(new_n306_), .C1(new_n563_), .C2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n278_), .A2(new_n215_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT35), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT74), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n221_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n278_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n608_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n600_), .A2(new_n605_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n607_), .B1(new_n617_), .B2(new_n610_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n612_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n615_), .B(KEYINPUT36), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n612_), .B2(new_n618_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT37), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n612_), .A2(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n620_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n612_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n273_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n212_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n212_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n631_), .B(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n636_), .B(KEYINPUT17), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n629_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n599_), .A2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT98), .Z(new_n647_));
  XOR2_X1   g446(.A(new_n513_), .B(KEYINPUT99), .Z(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n202_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n619_), .A2(new_n622_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT100), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n644_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n599_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n513_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n652_), .A2(new_n653_), .A3(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n560_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n203_), .B1(new_n658_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT39), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n647_), .A2(new_n203_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(new_n399_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n372_), .B1(new_n658_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT101), .Z(new_n671_));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n647_), .A2(new_n372_), .A3(new_n669_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n487_), .B(KEYINPUT102), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n658_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT42), .Z(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n677_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT103), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n647_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n654_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n644_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n599_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n513_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n306_), .A2(new_n233_), .A3(new_n686_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n629_), .B2(KEYINPUT104), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n563_), .A2(new_n598_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n629_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n629_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n697_), .B(new_n693_), .C1(new_n563_), .C2(new_n598_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n691_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n586_), .A2(new_n593_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n487_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n595_), .A2(new_n596_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n706_), .A2(new_n399_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n693_), .B1(new_n707_), .B2(new_n697_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n629_), .A3(new_n694_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n710_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n691_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n691_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n701_), .A2(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n649_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n690_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n688_), .A2(new_n717_), .A3(new_n662_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT45), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n701_), .A2(new_n711_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n560_), .B1(new_n713_), .B2(new_n712_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n723_), .B2(G36gat), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT106), .B(new_n717_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n719_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT46), .B(new_n719_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NAND3_X1  g529(.A1(new_n714_), .A2(G43gat), .A3(new_n669_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G43gat), .B1(new_n688_), .B2(new_n669_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g534(.A(G50gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n688_), .A2(new_n736_), .A3(new_n678_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n703_), .B1(new_n713_), .B2(new_n712_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n721_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n721_), .B2(new_n739_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n737_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT108), .B(new_n737_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1331gat));
  INV_X1    g546(.A(new_n306_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n707_), .A2(new_n232_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n657_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT109), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n752_), .A3(new_n657_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G57gat), .B1(new_n755_), .B2(new_n513_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n749_), .A2(new_n645_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n649_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1332gat));
  INV_X1    g559(.A(G64gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n761_), .A3(new_n662_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n751_), .A2(new_n662_), .A3(new_n753_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G64gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G64gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT110), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n757_), .A2(new_n769_), .A3(new_n669_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G71gat), .B1(new_n755_), .B2(new_n399_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT49), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT49), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(G1334gat));
  INV_X1    g573(.A(G78gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n757_), .A2(new_n775_), .A3(new_n678_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n678_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G78gat), .B1(new_n755_), .B2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(KEYINPUT50), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(KEYINPUT50), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  AND2_X1   g580(.A1(new_n749_), .A2(new_n687_), .ZN(new_n782_));
  INV_X1    g581(.A(G85gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n649_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n306_), .A2(new_n233_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n686_), .B(new_n785_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n689_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n787_), .B2(new_n783_), .ZN(G1336gat));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n662_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n560_), .A2(G92gat), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n789_), .A2(G92gat), .B1(new_n782_), .B2(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT111), .Z(G1337gat));
  NAND2_X1  g591(.A1(new_n786_), .A2(new_n669_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n669_), .A2(new_n251_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n793_), .A2(G99gat), .B1(new_n782_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n782_), .A2(new_n252_), .A3(new_n487_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n786_), .A2(new_n487_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(G106gat), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G106gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g603(.A(G113gat), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n233_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n212_), .A2(new_n216_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n211_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n210_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n210_), .A2(new_n809_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n609_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n222_), .B(KEYINPUT117), .C1(new_n216_), .C2(new_n212_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n219_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n230_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n231_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n820_), .A2(new_n302_), .A3(KEYINPUT119), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT119), .B1(new_n820_), .B2(new_n302_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n286_), .A2(new_n293_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n282_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n284_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(KEYINPUT55), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n300_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n301_), .A2(new_n232_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n301_), .B2(new_n232_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n829_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n654_), .B1(new_n823_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT57), .B1(new_n840_), .B2(KEYINPUT120), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n831_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n820_), .A2(new_n302_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n820_), .A2(new_n302_), .A3(KEYINPUT119), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n685_), .B1(new_n842_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n830_), .A2(KEYINPUT56), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n829_), .A2(new_n836_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n852_), .A2(new_n301_), .A3(new_n820_), .A4(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n697_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n855_), .B2(new_n854_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n841_), .A2(new_n851_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n644_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n232_), .A2(new_n644_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT114), .Z(new_n861_));
  NAND3_X1  g660(.A1(new_n748_), .A2(new_n861_), .A3(new_n697_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT54), .Z(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n648_), .B1(new_n859_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n560_), .A2(new_n488_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n863_), .B1(new_n858_), .B2(new_n644_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n866_), .A4(new_n648_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n806_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n859_), .A2(new_n864_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n867_), .A3(new_n649_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n873_), .B(new_n805_), .C1(new_n875_), .C2(new_n233_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n869_), .A2(new_n233_), .A3(new_n866_), .A4(new_n648_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT121), .B1(new_n877_), .B2(G113gat), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n872_), .A2(new_n876_), .A3(new_n878_), .ZN(G1340gat));
  NOR3_X1   g678(.A1(new_n869_), .A2(new_n866_), .A3(new_n648_), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n748_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n880_), .B(new_n882_), .C1(KEYINPUT60), .C2(new_n881_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n875_), .A2(new_n870_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n880_), .A2(KEYINPUT59), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n748_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n886_), .B2(new_n881_), .ZN(G1341gat));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n880_), .A2(new_n888_), .A3(new_n686_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n644_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n888_), .ZN(G1342gat));
  AOI21_X1  g690(.A(G134gat), .B1(new_n880_), .B2(new_n656_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n884_), .A2(new_n885_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(G134gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(G134gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n697_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n892_), .B1(new_n893_), .B2(new_n897_), .ZN(G1343gat));
  NOR3_X1   g697(.A1(new_n662_), .A2(new_n669_), .A3(new_n703_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n865_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n233_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n418_), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n748_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n419_), .ZN(G1345gat));
  NOR2_X1   g703(.A1(new_n900_), .A2(new_n644_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT61), .B(G155gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  NAND2_X1  g706(.A1(new_n629_), .A2(G162gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT123), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n865_), .A2(new_n899_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n899_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n869_), .A2(new_n648_), .A3(new_n655_), .A4(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(G162gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT124), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n910_), .B(new_n915_), .C1(new_n912_), .C2(G162gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1347gat));
  NOR3_X1   g716(.A1(new_n649_), .A2(new_n399_), .A3(new_n560_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(new_n777_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n874_), .A2(new_n232_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT22), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n925_));
  INV_X1    g724(.A(G169gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n920_), .B2(new_n924_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n923_), .B1(new_n925_), .B2(new_n927_), .ZN(G1348gat));
  NAND2_X1  g727(.A1(new_n874_), .A2(new_n919_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G176gat), .B1(new_n930_), .B2(new_n306_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n874_), .A2(KEYINPUT125), .A3(new_n703_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n869_), .B2(new_n487_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n932_), .A2(new_n918_), .A3(new_n934_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n306_), .A2(G176gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n931_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  NOR3_X1   g736(.A1(new_n929_), .A2(new_n521_), .A3(new_n644_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n932_), .A2(new_n934_), .A3(new_n686_), .A4(new_n918_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n349_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n929_), .B2(new_n697_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n656_), .A2(new_n383_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n929_), .B2(new_n942_), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n560_), .A2(new_n595_), .A3(new_n669_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n874_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n233_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n449_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n748_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n448_), .ZN(G1353gat));
  INV_X1    g748(.A(new_n945_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n644_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT126), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n954_), .B(KEYINPUT127), .Z(new_n955_));
  XNOR2_X1  g754(.A(new_n953_), .B(new_n955_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n945_), .B2(new_n697_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n656_), .A2(new_n456_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n945_), .B2(new_n958_), .ZN(G1355gat));
endmodule


