//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(G120gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT77), .ZN(new_n204_));
  INV_X1    g003(.A(G113gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(KEYINPUT77), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n202_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G113gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G120gat), .A3(new_n207_), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n217_), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  INV_X1    g017(.A(G155gat), .ZN(new_n219_));
  INV_X1    g018(.A(G162gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT80), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n216_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT81), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(new_n216_), .C1(new_n218_), .C2(new_n221_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT79), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G141gat), .ZN(new_n233_));
  INV_X1    g032(.A(G148gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n227_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n218_), .A2(new_n221_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(new_n228_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT83), .B(KEYINPUT2), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n232_), .B2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n235_), .B(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n238_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n215_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n237_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n214_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT98), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n210_), .A2(new_n213_), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n227_), .A2(new_n236_), .B1(new_n246_), .B2(new_n215_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n249_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n250_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT99), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G85gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  OR3_X1    g062(.A1(new_n257_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n249_), .A2(KEYINPUT4), .A3(new_n253_), .ZN(new_n265_));
  OR3_X1    g064(.A1(new_n251_), .A2(KEYINPUT4), .A3(new_n252_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n256_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n258_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT95), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT76), .B(G176gat), .ZN(new_n271_));
  INV_X1    g070(.A(G169gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT22), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G169gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT93), .B1(new_n273_), .B2(new_n275_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n271_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT94), .ZN(new_n287_));
  INV_X1    g086(.A(new_n285_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(new_n282_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n284_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n280_), .A2(new_n281_), .A3(new_n287_), .A4(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n296_));
  OAI22_X1  g095(.A1(new_n293_), .A2(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT92), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT92), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n289_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n281_), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n302_), .B(new_n305_), .C1(new_n299_), .C2(new_n301_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n292_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G197gat), .ZN(new_n311_));
  INV_X1    g110(.A(G197gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G204gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(G211gat), .A2(G218gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G211gat), .A2(G218gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT87), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G211gat), .ZN(new_n318_));
  INV_X1    g117(.A(G218gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G211gat), .A2(G218gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT88), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n323_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n311_), .A2(new_n313_), .A3(new_n309_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n311_), .A2(new_n313_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT21), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n314_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT88), .A3(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n270_), .B1(new_n308_), .B2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n332_), .A2(new_n327_), .B1(new_n324_), .B2(KEYINPUT88), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n330_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n304_), .A2(new_n306_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n276_), .A2(new_n277_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT93), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n305_), .B1(new_n344_), .B2(new_n271_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n287_), .A2(new_n291_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n340_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n339_), .A2(new_n347_), .A3(KEYINPUT95), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  INV_X1    g148(.A(new_n302_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(KEYINPUT24), .A3(new_n281_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n302_), .A2(new_n298_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n297_), .A2(new_n289_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n271_), .B1(new_n342_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n354_), .B2(new_n273_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n286_), .A2(new_n281_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n349_), .B1(new_n334_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n335_), .A2(new_n348_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n334_), .A2(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n308_), .A2(new_n334_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT20), .A4(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G64gat), .ZN(new_n371_));
  INV_X1    g170(.A(G92gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT96), .ZN(new_n375_));
  INV_X1    g174(.A(new_n373_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n364_), .A2(new_n376_), .A3(new_n367_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n368_), .A2(KEYINPUT96), .A3(new_n373_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n265_), .A2(G225gat), .A3(G233gat), .A4(new_n266_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n249_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n263_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT33), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n269_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n331_), .A2(new_n386_), .A3(new_n333_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n248_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n252_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n395_), .B(KEYINPUT85), .Z(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n392_), .B1(new_n237_), .B2(new_n247_), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n396_), .B(KEYINPUT86), .Z(new_n399_));
  NOR3_X1   g198(.A1(new_n398_), .A2(new_n339_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n397_), .A2(new_n403_), .A3(new_n401_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT91), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n403_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n409_));
  AOI211_X1 g208(.A(new_n404_), .B(new_n400_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n252_), .A2(new_n392_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G22gat), .B(G50gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n413_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n407_), .A2(new_n411_), .A3(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n421_), .B(new_n408_), .C1(new_n410_), .C2(new_n409_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n381_), .A2(new_n382_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n263_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT100), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n383_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n381_), .A2(KEYINPUT100), .A3(new_n263_), .A4(new_n382_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n368_), .B1(new_n431_), .B2(new_n376_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n365_), .A2(KEYINPUT20), .A3(new_n366_), .A4(new_n363_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n347_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n434_), .A2(new_n359_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n363_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT32), .A3(new_n373_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .A4(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n385_), .A2(new_n425_), .A3(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n423_), .A2(new_n424_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n429_), .A2(new_n430_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n378_), .A2(new_n442_), .A3(new_n379_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n376_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n440_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n358_), .B(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT30), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G15gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n450_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n448_), .B(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(KEYINPUT78), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(KEYINPUT78), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n214_), .B(KEYINPUT31), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n456_), .A2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n439_), .A2(new_n447_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n429_), .A2(new_n430_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n443_), .A2(new_n445_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n466_), .A2(KEYINPUT101), .A3(new_n425_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT101), .B1(new_n466_), .B2(new_n425_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n465_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT102), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT101), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(KEYINPUT101), .A3(new_n425_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(KEYINPUT102), .A3(new_n465_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n461_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT65), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n482_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT7), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G85gat), .B(G92gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n478_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT66), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n485_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n478_), .A3(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(KEYINPUT66), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT9), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(G85gat), .A3(G92gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT10), .B(G99gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(G106gat), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n501_), .A2(new_n503_), .A3(new_n483_), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n504_), .B(KEYINPUT64), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n509_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n498_), .A2(new_n505_), .A3(new_n513_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n513_), .B(KEYINPUT67), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n506_), .A2(KEYINPUT12), .A3(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n518_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n519_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n513_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n522_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n539_), .B2(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT71), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G29gat), .B(G36gat), .ZN(new_n546_));
  INV_X1    g345(.A(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G50gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT15), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G1gat), .B(G8gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT72), .ZN(new_n553_));
  INV_X1    g352(.A(G15gat), .ZN(new_n554_));
  INV_X1    g353(.A(G22gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G15gat), .A2(G22gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G1gat), .A2(G8gat), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n556_), .A2(new_n557_), .B1(KEYINPUT14), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n553_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n551_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n550_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT74), .Z(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n560_), .B(new_n550_), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(G229gat), .A3(G233gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n272_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n312_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n477_), .A2(new_n545_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n506_), .A2(new_n551_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  OAI221_X1 g381(.A(new_n580_), .B1(KEYINPUT35), .B2(new_n582_), .C1(new_n562_), .C2(new_n506_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G134gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n220_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n590_), .B(new_n591_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n594_), .A3(new_n586_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n579_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(new_n579_), .A3(new_n595_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n560_), .B(new_n600_), .Z(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(new_n520_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n520_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G183gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n318_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n602_), .A2(new_n603_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n601_), .B(new_n513_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT73), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n599_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n578_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT103), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n620_), .A2(G1gat), .A3(new_n462_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n622_));
  INV_X1    g421(.A(new_n545_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n439_), .A2(new_n447_), .A3(new_n460_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT102), .B1(new_n475_), .B2(new_n465_), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n470_), .B(new_n464_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n627_), .A3(new_n576_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n593_), .A2(new_n595_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n628_), .A2(new_n617_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n462_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n622_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(G8gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n630_), .B2(new_n446_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT39), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n620_), .A2(G8gat), .A3(new_n466_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1325gat));
  AOI21_X1  g441(.A(new_n554_), .B1(new_n630_), .B2(new_n463_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n628_), .A2(new_n617_), .A3(new_n599_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n554_), .A3(new_n463_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1326gat));
  AOI21_X1  g446(.A(new_n555_), .B1(new_n630_), .B2(new_n440_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT42), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n555_), .A3(new_n440_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1327gat));
  INV_X1    g450(.A(new_n629_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n616_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n578_), .A2(new_n653_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n654_), .A2(G29gat), .A3(new_n462_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n542_), .A2(new_n576_), .A3(new_n544_), .A4(new_n617_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n599_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n598_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n596_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n477_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n662_), .B2(KEYINPUT104), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n627_), .B2(new_n599_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n657_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n660_), .B1(new_n477_), .B2(new_n662_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n627_), .A2(new_n599_), .A3(new_n664_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n656_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT44), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n441_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(G29gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n673_), .B2(G29gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n655_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g477(.A(new_n654_), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n446_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n667_), .B(new_n656_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n466_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n680_), .B1(new_n686_), .B2(new_n668_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n683_), .A2(new_n684_), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n683_), .B2(new_n687_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  NAND4_X1  g489(.A1(new_n668_), .A2(G43gat), .A3(new_n672_), .A4(new_n463_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n547_), .B1(new_n654_), .B2(new_n460_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n691_), .A2(new_n692_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT107), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT47), .B1(new_n700_), .B2(new_n694_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1330gat));
  NAND3_X1  g501(.A1(new_n679_), .A2(new_n549_), .A3(new_n440_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n668_), .A2(new_n440_), .A3(new_n672_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G50gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n440_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n704_), .B(G50gat), .C1(new_n707_), .C2(new_n685_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n703_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n712_), .B(new_n703_), .C1(new_n706_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1331gat));
  NOR3_X1   g513(.A1(new_n623_), .A2(new_n477_), .A3(new_n576_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n629_), .A2(new_n617_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(G57gat), .A3(new_n441_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT110), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n715_), .A2(new_n618_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n441_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n723_), .A3(new_n446_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n717_), .A2(new_n446_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G64gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT48), .B(new_n723_), .C1(new_n717_), .C2(new_n446_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(G1333gat));
  NOR2_X1   g529(.A1(new_n460_), .A2(G71gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT112), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n720_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n717_), .A2(new_n463_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G71gat), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT49), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT49), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n720_), .A2(new_n739_), .A3(new_n440_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n717_), .A2(new_n440_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G78gat), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT50), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT50), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  AND2_X1   g544(.A1(new_n715_), .A2(new_n653_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n441_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n669_), .A2(new_n670_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n623_), .A2(new_n576_), .A3(new_n616_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n441_), .A2(G85gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n747_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  AOI21_X1  g553(.A(G92gat), .B1(new_n746_), .B2(new_n446_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n466_), .A2(new_n372_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n752_), .B2(new_n756_), .ZN(G1337gat));
  NAND4_X1  g556(.A1(new_n749_), .A2(new_n463_), .A3(new_n750_), .A4(new_n751_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G99gat), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n460_), .A2(new_n502_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT114), .B1(new_n746_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g562(.A(G106gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n764_), .A3(new_n440_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n748_), .A2(new_n750_), .A3(new_n440_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n519_), .B1(new_n525_), .B2(KEYINPUT12), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n506_), .A2(KEYINPUT12), .A3(new_n520_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n523_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n774_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n523_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n774_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n522_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n532_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n534_), .A2(new_n577_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n786_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n532_), .B(new_n789_), .C1(new_n780_), .C2(new_n783_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n787_), .A2(KEYINPUT117), .A3(new_n788_), .A4(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n567_), .A2(new_n565_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n561_), .A2(new_n563_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n565_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n575_), .B1(new_n797_), .B2(new_n574_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT118), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n536_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n793_), .A2(new_n794_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n652_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n784_), .A2(KEYINPUT56), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n534_), .B1(new_n784_), .B2(KEYINPUT56), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n799_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT58), .A4(new_n799_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n599_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n801_), .A2(KEYINPUT57), .A3(new_n652_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n662_), .A2(new_n577_), .A3(new_n616_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n541_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OR3_X1    g615(.A1(new_n814_), .A2(KEYINPUT54), .A3(new_n815_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n813_), .A2(new_n617_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n475_), .A2(new_n441_), .A3(new_n463_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT119), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n576_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n818_), .A2(KEYINPUT120), .A3(new_n825_), .A4(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT121), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n817_), .A2(new_n816_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n812_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT57), .B1(new_n801_), .B2(new_n652_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n811_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n616_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n820_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n825_), .B1(new_n835_), .B2(KEYINPUT120), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n821_), .A2(new_n823_), .A3(KEYINPUT59), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n827_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n576_), .A2(KEYINPUT122), .A3(G113gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(KEYINPUT122), .B2(G113gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n822_), .B1(new_n840_), .B2(new_n842_), .ZN(G1340gat));
  XOR2_X1   g642(.A(KEYINPUT123), .B(G120gat), .Z(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n623_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n821_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n623_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n821_), .B2(new_n616_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n616_), .A2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n840_), .B2(new_n850_), .ZN(G1342gat));
  AOI21_X1  g650(.A(G134gat), .B1(new_n821_), .B2(new_n629_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n599_), .A2(G134gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n840_), .B2(new_n853_), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n818_), .A2(new_n463_), .A3(new_n425_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n462_), .A2(new_n446_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n577_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n233_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n623_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n234_), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n857_), .A2(new_n617_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT124), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n862_), .B(new_n864_), .ZN(G1346gat));
  NOR3_X1   g664(.A1(new_n857_), .A2(new_n220_), .A3(new_n662_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n857_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n629_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n220_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n441_), .A2(new_n466_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n440_), .A2(new_n460_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n833_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n872_), .A2(new_n576_), .A3(new_n344_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n272_), .B1(new_n872_), .B2(new_n576_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT62), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(KEYINPUT62), .B2(new_n874_), .ZN(G1348gat));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n545_), .ZN(new_n877_));
  INV_X1    g676(.A(G176gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n271_), .B2(new_n877_), .ZN(G1349gat));
  INV_X1    g679(.A(new_n872_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G183gat), .B1(new_n881_), .B2(new_n617_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n872_), .B(new_n616_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1350gat));
  OAI211_X1 g683(.A(new_n872_), .B(new_n629_), .C1(new_n296_), .C2(new_n295_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n872_), .A2(new_n599_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n886_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT125), .B1(new_n886_), .B2(G190gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n885_), .B1(new_n887_), .B2(new_n888_), .ZN(G1351gat));
  NAND4_X1  g688(.A1(new_n833_), .A2(new_n460_), .A3(new_n440_), .A4(new_n870_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n818_), .A2(new_n425_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n460_), .A4(new_n870_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G197gat), .B1(new_n895_), .B2(new_n576_), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n312_), .B(new_n577_), .C1(new_n891_), .C2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1352gat));
  AOI21_X1  g697(.A(new_n893_), .B1(new_n855_), .B2(new_n870_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n545_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G204gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n895_), .A2(new_n310_), .A3(new_n545_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1353gat));
  OR2_X1    g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n895_), .B2(new_n616_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n617_), .B(new_n907_), .C1(new_n891_), .C2(new_n894_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1354gat));
  XOR2_X1   g708(.A(KEYINPUT127), .B(G218gat), .Z(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n895_), .B2(new_n629_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n910_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n662_), .B(new_n912_), .C1(new_n891_), .C2(new_n894_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1355gat));
endmodule


