//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  INV_X1    g014(.A(new_n208_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT82), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n215_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n222_), .A3(KEYINPUT83), .A4(KEYINPUT24), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n214_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT79), .B(G183gat), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT25), .ZN(new_n229_));
  INV_X1    g028(.A(G190gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT80), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT26), .ZN(new_n232_));
  INV_X1    g031(.A(G183gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n229_), .B(new_n232_), .C1(KEYINPUT25), .C2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n206_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n222_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n213_), .B1(G190gat), .B2(new_n227_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n226_), .A2(new_n234_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242_));
  INV_X1    g041(.A(G197gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(G204gat), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G197gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT21), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT87), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n245_), .A3(G197gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT87), .B1(new_n243_), .B2(G204gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(new_n244_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n242_), .B(new_n247_), .C1(new_n251_), .C2(KEYINPUT21), .ZN(new_n252_));
  INV_X1    g051(.A(new_n242_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT21), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n203_), .B1(new_n241_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n257_));
  INV_X1    g056(.A(new_n255_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n259_), .A2(new_n213_), .A3(new_n211_), .A4(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n211_), .A2(new_n213_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(KEYINPUT89), .A3(new_n259_), .A4(new_n262_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n233_), .A2(new_n230_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n213_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(new_n237_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n257_), .B(new_n258_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT90), .B1(new_n273_), .B2(new_n255_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n256_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT19), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT88), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  AOI211_X1 g078(.A(new_n203_), .B(new_n277_), .C1(new_n273_), .C2(new_n255_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n226_), .A2(new_n234_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n239_), .A2(new_n240_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n258_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287_));
  INV_X1    g086(.A(G92gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT18), .B(G64gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT32), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n202_), .B1(new_n286_), .B2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n255_), .B(new_n263_), .C1(new_n237_), .C2(new_n270_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT20), .B(new_n296_), .C1(new_n241_), .C2(new_n255_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n277_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  OR2_X1    g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n300_), .B(new_n301_), .C1(new_n304_), .C2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n302_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n301_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n309_), .B(new_n305_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315_));
  XOR2_X1   g114(.A(G113gat), .B(G120gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n314_), .B(new_n318_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n319_), .B(new_n321_), .C1(new_n322_), .C2(new_n315_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G57gat), .B(G85gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n324_), .A3(new_n332_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n299_), .A2(new_n294_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n275_), .A2(new_n278_), .B1(new_n284_), .B2(new_n280_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT96), .A3(new_n293_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n295_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT97), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n295_), .A2(KEYINPUT97), .A3(new_n334_), .A4(new_n336_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n319_), .B(new_n320_), .C1(new_n322_), .C2(new_n315_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n320_), .B1(new_n322_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n344_), .B2(new_n322_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n330_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT33), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n347_), .A2(KEYINPUT95), .B1(new_n348_), .B2(new_n333_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n333_), .A2(new_n348_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT91), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n335_), .B2(new_n292_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n279_), .A2(new_n292_), .A3(new_n285_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n286_), .A2(new_n351_), .A3(new_n291_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n349_), .B(new_n350_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n347_), .A2(KEYINPUT95), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n339_), .B(new_n340_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G22gat), .B(G50gat), .Z(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n255_), .B1(KEYINPUT29), .B2(new_n314_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n314_), .A2(KEYINPUT29), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n367_), .A2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n364_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n369_), .A3(new_n363_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n318_), .B(KEYINPUT31), .Z(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(G15gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G43gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(G71gat), .B(G99gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n283_), .A2(KEYINPUT30), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n241_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n383_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n383_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n376_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n387_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n241_), .A2(new_n386_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT85), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n382_), .B1(new_n397_), .B2(new_n388_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n376_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n398_), .A2(new_n392_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n375_), .B1(new_n394_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n353_), .A2(KEYINPUT98), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n299_), .B2(new_n291_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT98), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n354_), .A2(new_n355_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n404_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n331_), .A2(new_n333_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n372_), .A2(new_n374_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n399_), .B1(new_n398_), .B2(new_n392_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n391_), .A2(new_n393_), .A3(new_n376_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n401_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n358_), .A2(new_n402_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G230gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT64), .ZN(new_n420_));
  INV_X1    g219(.A(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(G99gat), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(KEYINPUT10), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(KEYINPUT10), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G85gat), .A2(G92gat), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n426_), .A2(KEYINPUT9), .ZN(new_n427_));
  INV_X1    g226(.A(G85gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n288_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(KEYINPUT9), .A3(new_n426_), .ZN(new_n430_));
  AND3_X1   g229(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n425_), .A2(new_n427_), .A3(new_n430_), .A4(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT7), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(new_n422_), .A3(new_n421_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G99gat), .A2(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n436_), .A2(new_n439_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT8), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n429_), .A2(new_n426_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n434_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n448_));
  INV_X1    g247(.A(G57gat), .ZN(new_n449_));
  INV_X1    g248(.A(G64gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G57gat), .A2(G64gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G71gat), .B(G78gat), .Z(new_n454_));
  OR2_X1    g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n451_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n456_), .B2(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n420_), .B1(new_n447_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT65), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n442_), .A2(new_n444_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n433_), .A2(new_n430_), .A3(new_n427_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n463_), .A2(new_n464_), .B1(new_n425_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n458_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n461_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n447_), .A2(KEYINPUT12), .A3(new_n458_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT65), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n470_), .B(new_n420_), .C1(new_n447_), .C2(new_n458_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n460_), .A2(new_n468_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n420_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n467_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n466_), .A2(new_n467_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT5), .B(G176gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G204gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G120gat), .B(G148gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n472_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n472_), .A2(KEYINPUT66), .A3(new_n477_), .A4(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT13), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(KEYINPUT67), .A3(new_n488_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n486_), .B2(new_n488_), .ZN(new_n495_));
  AOI211_X1 g294(.A(new_n490_), .B(new_n487_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT13), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G29gat), .B(G36gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n500_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT78), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508_));
  INV_X1    g307(.A(G1gat), .ZN(new_n509_));
  INV_X1    g308(.A(G8gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G1gat), .B(G8gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n506_), .B(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n514_), .ZN(new_n519_));
  OAI211_X1 g318(.A(G229gat), .B(G233gat), .C1(new_n516_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n514_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n506_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n515_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n520_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n520_), .B2(new_n526_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n499_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n418_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G127gat), .B(G155gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G211gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT16), .B(G183gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT77), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n458_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n458_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n546_));
  OAI211_X1 g345(.A(G231gat), .B(G233gat), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n514_), .B(KEYINPUT76), .ZN(new_n548_));
  INV_X1    g347(.A(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n544_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT73), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT71), .B(KEYINPUT72), .Z(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT74), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n447_), .A2(KEYINPUT69), .A3(new_n506_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n523_), .A2(new_n447_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT69), .B1(new_n447_), .B2(new_n506_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT34), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(KEYINPUT35), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(KEYINPUT35), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n572_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581_));
  INV_X1    g380(.A(new_n576_), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n581_), .B(new_n582_), .C1(new_n570_), .C2(new_n573_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n572_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n568_), .B1(new_n580_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n583_), .B2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n577_), .A2(new_n572_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n563_), .A2(new_n564_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n587_), .A2(new_n588_), .A3(new_n566_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT75), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n594_), .A3(KEYINPUT37), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n586_), .B(new_n591_), .C1(new_n593_), .C2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n555_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n537_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n509_), .A3(new_n411_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT38), .ZN(new_n602_));
  INV_X1    g401(.A(new_n592_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n555_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n537_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n412_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(G1324gat));
  INV_X1    g406(.A(new_n605_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n410_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G8gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n600_), .A2(new_n510_), .A3(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n610_), .A2(G8gat), .A3(new_n616_), .A4(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT40), .Z(G1325gat));
  NOR2_X1   g419(.A1(new_n400_), .A2(new_n394_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G15gat), .B1(new_n605_), .B2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT41), .Z(new_n624_));
  NAND3_X1  g423(.A1(new_n600_), .A2(new_n378_), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n600_), .A2(new_n627_), .A3(new_n413_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n608_), .B2(new_n413_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n629_), .A2(new_n630_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT100), .Z(G1327gat));
  INV_X1    g434(.A(new_n555_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n595_), .A2(new_n597_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT43), .B1(new_n418_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n339_), .A2(new_n340_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n352_), .B(new_n353_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n357_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n350_), .A4(new_n349_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n401_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n642_), .A2(KEYINPUT27), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n401_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n408_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n640_), .B(new_n637_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n536_), .B(new_n636_), .C1(new_n639_), .C2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT101), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n639_), .A2(new_n649_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n535_), .A3(new_n555_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n650_), .A2(KEYINPUT44), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n657_), .A2(new_n411_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(G29gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n603_), .A2(new_n555_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT102), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n537_), .A2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n411_), .A2(new_n660_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT104), .Z(new_n669_));
  OAI22_X1  g468(.A1(new_n659_), .A2(new_n660_), .B1(new_n667_), .B2(new_n669_), .ZN(G1328gat));
  XNOR2_X1  g469(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n410_), .B1(new_n651_), .B2(new_n656_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n658_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n665_), .A2(new_n673_), .A3(new_n666_), .A4(new_n609_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n656_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n654_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n609_), .B(new_n658_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n671_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n685_), .ZN(G1329gat));
  NAND4_X1  g485(.A1(new_n657_), .A2(G43gat), .A3(new_n621_), .A4(new_n658_), .ZN(new_n687_));
  INV_X1    g486(.A(G43gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(new_n667_), .B2(new_n622_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT47), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1330gat));
  NOR2_X1   g493(.A1(new_n375_), .A2(G50gat), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT107), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n665_), .A2(new_n666_), .A3(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n657_), .A2(new_n413_), .A3(new_n658_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1331gat));
  NAND2_X1  g501(.A1(new_n358_), .A2(new_n402_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n609_), .B2(new_n647_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n534_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT108), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(new_n499_), .A3(new_n598_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n449_), .A3(new_n411_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n534_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n498_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n704_), .A2(new_n604_), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n412_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1332gat));
  OAI21_X1  g514(.A(G64gat), .B1(new_n711_), .B2(new_n410_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT48), .ZN(new_n717_));
  INV_X1    g516(.A(new_n707_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n609_), .A2(new_n450_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n711_), .B2(new_n622_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT49), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n622_), .A2(G71gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n718_), .B2(new_n723_), .ZN(G1334gat));
  OAI21_X1  g523(.A(G78gat), .B1(new_n711_), .B2(new_n375_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT50), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n375_), .A2(G78gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n718_), .B2(new_n727_), .ZN(G1335gat));
  NAND3_X1  g527(.A1(new_n706_), .A2(new_n499_), .A3(new_n663_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(new_n412_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n652_), .A2(new_n555_), .A3(new_n710_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n411_), .A2(G85gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT110), .Z(new_n733_));
  AOI22_X1  g532(.A1(new_n730_), .A2(new_n428_), .B1(new_n731_), .B2(new_n733_), .ZN(G1336gat));
  OAI21_X1  g533(.A(new_n288_), .B1(new_n729_), .B2(new_n410_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n735_), .A2(KEYINPUT111), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(KEYINPUT111), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n410_), .A2(new_n288_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n736_), .A2(new_n737_), .B1(new_n731_), .B2(new_n738_), .ZN(G1337gat));
  NAND2_X1  g538(.A1(new_n731_), .A2(new_n621_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT112), .B1(new_n740_), .B2(G99gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n621_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n741_), .A2(new_n742_), .B1(new_n729_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  OAI221_X1 g546(.A(new_n745_), .B1(new_n729_), .B2(new_n743_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1338gat));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n731_), .A2(new_n413_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G106gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT52), .B(new_n421_), .C1(new_n731_), .C2(new_n413_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n413_), .A2(new_n421_), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n752_), .A2(new_n753_), .B1(new_n729_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT53), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757_));
  OAI221_X1 g556(.A(new_n757_), .B1(new_n729_), .B2(new_n754_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n709_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n598_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(new_n598_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n498_), .A2(new_n598_), .A3(new_n534_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n761_), .A2(new_n762_), .A3(new_n598_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(KEYINPUT54), .A3(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n765_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n534_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n468_), .A2(new_n474_), .A3(new_n469_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n473_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(new_n473_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n472_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n472_), .A2(KEYINPUT115), .A3(new_n777_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n472_), .A2(new_n777_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n776_), .A2(new_n780_), .A3(new_n781_), .A4(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n481_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n784_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n771_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT117), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n525_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n521_), .A2(new_n524_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n789_), .B(new_n529_), .C1(new_n525_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n531_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n771_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n788_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n785_), .A2(new_n786_), .A3(KEYINPUT118), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n783_), .A2(new_n784_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(KEYINPUT118), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n486_), .A3(new_n793_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n786_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n784_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n792_), .B1(new_n786_), .B2(KEYINPUT118), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(KEYINPUT58), .A4(new_n486_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n805_), .A2(new_n637_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n797_), .B2(new_n592_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n798_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n770_), .B1(new_n814_), .B2(new_n636_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n609_), .A2(new_n412_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n621_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n819_));
  NAND4_X1  g618(.A1(new_n815_), .A2(new_n375_), .A3(new_n818_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n765_), .A2(new_n769_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n797_), .A2(new_n592_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n805_), .A2(new_n637_), .A3(new_n811_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n821_), .B1(new_n827_), .B2(new_n555_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n828_), .A2(new_n413_), .A3(new_n817_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(KEYINPUT59), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n820_), .B(new_n709_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G113gat), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n834_), .A3(new_n709_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT120), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n838_), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n498_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n829_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n829_), .A2(new_n831_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n844_), .A2(new_n499_), .A3(new_n820_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n829_), .B2(new_n636_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n844_), .A2(new_n820_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n636_), .A2(G127gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT121), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n848_), .B2(new_n850_), .ZN(G1342gat));
  AND2_X1   g650(.A1(new_n829_), .A2(new_n603_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(G134gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n844_), .A2(G134gat), .A3(new_n637_), .A4(new_n820_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1343gat));
  NOR3_X1   g654(.A1(new_n828_), .A2(new_n621_), .A3(new_n375_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n816_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n709_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n857_), .A2(new_n498_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT122), .B(G148gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1345gat));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT123), .B1(new_n857_), .B2(new_n555_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n555_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n865_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n555_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n866_), .A3(new_n864_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1346gat));
  AND3_X1   g671(.A1(new_n858_), .A2(G162gat), .A3(new_n637_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G162gat), .B1(new_n858_), .B2(new_n603_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n828_), .A2(new_n413_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n410_), .A2(new_n411_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n876_), .A2(new_n621_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n709_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n621_), .A3(new_n877_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881_), .B2(new_n534_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n235_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n880_), .B(new_n884_), .C1(new_n885_), .C2(new_n879_), .ZN(G1348gat));
  OR2_X1    g685(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n878_), .A2(new_n499_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT125), .Z(new_n890_));
  XOR2_X1   g689(.A(new_n888_), .B(new_n890_), .Z(G1349gat));
  NOR2_X1   g690(.A1(new_n881_), .A2(new_n555_), .ZN(new_n892_));
  MUX2_X1   g691(.A(new_n227_), .B(new_n260_), .S(new_n892_), .Z(G1350gat));
  NAND3_X1  g692(.A1(new_n878_), .A2(new_n261_), .A3(new_n603_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G190gat), .B1(new_n881_), .B2(new_n638_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NAND3_X1  g695(.A1(new_n856_), .A2(new_n709_), .A3(new_n877_), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n897_), .A2(KEYINPUT126), .A3(new_n243_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n243_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT126), .B1(new_n897_), .B2(new_n243_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .ZN(G1352gat));
  AND2_X1   g700(.A1(new_n856_), .A2(new_n877_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n499_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT127), .B(G204gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1353gat));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n902_), .B(new_n636_), .C1(new_n906_), .C2(new_n907_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n902_), .A2(new_n636_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n906_), .ZN(G1354gat));
  AOI21_X1  g709(.A(G218gat), .B1(new_n902_), .B2(new_n603_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n902_), .A2(G218gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n637_), .B2(new_n912_), .ZN(G1355gat));
endmodule


