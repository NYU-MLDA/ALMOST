//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n203_), .B(new_n204_), .C1(new_n207_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n205_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(new_n204_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n212_), .B(new_n208_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT86), .ZN(new_n218_));
  XOR2_X1   g017(.A(G113gat), .B(G120gat), .Z(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n217_), .A2(new_n221_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n202_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT4), .B1(new_n218_), .B2(new_n221_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G225gat), .A2(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT94), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT94), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n222_), .A2(new_n223_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n227_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n236_));
  XNOR2_X1  g035(.A(G1gat), .B(G29gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G85gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n229_), .A2(new_n232_), .A3(new_n240_), .A4(new_n234_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT27), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT20), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n247_));
  XNOR2_X1  g046(.A(G197gat), .B(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT91), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(KEYINPUT91), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(KEYINPUT89), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G169gat), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT83), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n267_));
  OAI22_X1  g066(.A1(new_n265_), .A2(new_n266_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G183gat), .ZN(new_n269_));
  INV_X1    g068(.A(G190gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n263_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n274_));
  AND2_X1   g073(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G169gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n260_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT24), .A3(new_n262_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(KEYINPUT24), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n265_), .A2(new_n266_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n272_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n246_), .B1(new_n258_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT19), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n253_), .A2(new_n257_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n262_), .B(new_n261_), .C1(new_n282_), .C2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n268_), .A2(new_n279_), .A3(new_n280_), .A4(new_n276_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n289_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(new_n288_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT93), .ZN(new_n295_));
  XOR2_X1   g094(.A(G8gat), .B(G36gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G92gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT18), .B(G64gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n272_), .A2(new_n283_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n289_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n291_), .A2(new_n292_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n302_), .B(KEYINPUT20), .C1(new_n289_), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n287_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT93), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n285_), .A2(new_n306_), .A3(new_n288_), .A4(new_n293_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n295_), .A2(new_n300_), .A3(new_n305_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT96), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n285_), .A2(new_n293_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n287_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n287_), .B2(new_n304_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n299_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n245_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n295_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n299_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n317_), .A2(new_n308_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n318_), .A2(new_n245_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT97), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(G228gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(G228gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n289_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n326_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n217_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n329_), .B1(new_n334_), .B2(new_n289_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n218_), .A2(KEYINPUT29), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G78gat), .B(G106gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  AND2_X1   g143(.A1(new_n335_), .A2(new_n336_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n335_), .A2(new_n336_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n339_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n221_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT85), .B(G71gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT84), .B(G99gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G15gat), .B(G43gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT30), .B(KEYINPUT31), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n301_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n356_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n349_), .A2(new_n350_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT97), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n318_), .A2(new_n245_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n308_), .A2(KEYINPUT96), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n308_), .A2(KEYINPUT96), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n366_), .A2(new_n314_), .A3(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n364_), .B(new_n365_), .C1(new_n368_), .C2(new_n245_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n320_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n350_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n348_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n372_), .B(new_n362_), .C1(new_n315_), .C2(new_n319_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n244_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n300_), .A2(KEYINPUT32), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n313_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n244_), .B(new_n376_), .C1(new_n316_), .C2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n226_), .A2(new_n227_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n233_), .A2(new_n228_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n241_), .A3(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n243_), .A2(KEYINPUT33), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n243_), .A2(KEYINPUT33), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n318_), .B(new_n380_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  AOI211_X1 g182(.A(new_n361_), .B(new_n372_), .C1(new_n377_), .C2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n374_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G230gat), .A2(G233gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT64), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G71gat), .B(G78gat), .Z(new_n389_));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G57gat), .A2(G64gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G57gat), .A2(G64gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G57gat), .ZN(new_n395_));
  INV_X1    g194(.A(G64gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(KEYINPUT67), .A3(new_n391_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n394_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n389_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(new_n389_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT66), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT7), .ZN(new_n407_));
  INV_X1    g206(.A(G99gat), .ZN(new_n408_));
  INV_X1    g207(.A(G106gat), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .A4(KEYINPUT65), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n411_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n410_), .A2(new_n412_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(G85gat), .A2(G92gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G85gat), .A2(G92gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n406_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT8), .ZN(new_n422_));
  INV_X1    g221(.A(new_n416_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(KEYINPUT9), .A3(new_n419_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n419_), .A2(KEYINPUT9), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT10), .B(G99gat), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n409_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n421_), .A2(new_n422_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n417_), .A2(new_n420_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT66), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n410_), .A2(new_n412_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n415_), .A2(new_n416_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n406_), .B(new_n420_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(KEYINPUT8), .A3(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n405_), .A2(KEYINPUT68), .A3(new_n431_), .A4(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(KEYINPUT66), .A3(new_n422_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n428_), .A2(new_n430_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(KEYINPUT8), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n440_), .B(new_n441_), .C1(new_n442_), .C2(new_n421_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n443_), .B2(new_n404_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n438_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n404_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n388_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT69), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(new_n404_), .A3(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n431_), .A2(new_n437_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n388_), .B1(new_n443_), .B2(new_n404_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT5), .B(G176gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G204gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(G120gat), .B(G148gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  OR3_X1    g258(.A1(new_n447_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n447_), .B2(new_n455_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT13), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G29gat), .B(G36gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G43gat), .B(G50gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT80), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G1gat), .A2(G8gat), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n474_), .A2(KEYINPUT77), .A3(KEYINPUT14), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT77), .B1(new_n474_), .B2(KEYINPUT14), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n472_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT81), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n472_), .B2(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n471_), .B(KEYINPUT15), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n481_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n483_), .A2(new_n485_), .B1(new_n481_), .B2(new_n472_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(new_n487_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n490_), .B(new_n498_), .C1(new_n487_), .C2(new_n492_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n464_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n385_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n404_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n481_), .B(KEYINPUT78), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G183gat), .B(G211gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(G127gat), .B(G155gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT17), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n514_), .A2(KEYINPUT17), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n509_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n515_), .B2(new_n509_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n443_), .A2(new_n471_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT34), .Z(new_n522_));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT71), .Z(new_n525_));
  AND2_X1   g324(.A1(new_n520_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n488_), .A2(new_n443_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(new_n523_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT73), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n520_), .A2(new_n527_), .A3(new_n525_), .A4(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n488_), .A2(new_n531_), .A3(new_n443_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(KEYINPUT70), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n526_), .A2(new_n530_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n536_));
  XOR2_X1   g335(.A(G134gat), .B(G162gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(G218gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT72), .B(G190gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n530_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n535_), .A2(new_n536_), .A3(new_n540_), .A4(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n534_), .B2(new_n528_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n540_), .B(KEYINPUT36), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT74), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n544_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n543_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT75), .B1(new_n535_), .B2(new_n543_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n547_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT76), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n556_), .B(new_n547_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n544_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n551_), .B1(new_n558_), .B2(new_n550_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n505_), .A2(new_n519_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n244_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n560_), .A2(G1gat), .A3(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT38), .Z(new_n563_));
  OR2_X1    g362(.A1(new_n374_), .A2(new_n384_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n564_), .A2(new_n519_), .A3(new_n503_), .A4(new_n558_), .ZN(new_n565_));
  OAI21_X1  g364(.A(G1gat), .B1(new_n565_), .B2(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(G1324gat));
  INV_X1    g366(.A(KEYINPUT39), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n320_), .A2(new_n369_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n568_), .B(G8gat), .C1(new_n565_), .C2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT99), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n503_), .B(new_n558_), .C1(new_n374_), .C2(new_n384_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n574_), .A2(new_n518_), .A3(new_n570_), .ZN(new_n575_));
  INV_X1    g374(.A(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT39), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT98), .B(KEYINPUT39), .C1(new_n575_), .C2(new_n576_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n575_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n581_), .A2(KEYINPUT99), .A3(new_n568_), .A4(G8gat), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n573_), .A2(new_n579_), .A3(new_n580_), .A4(new_n582_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n560_), .A2(G8gat), .A3(new_n570_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(KEYINPUT40), .A3(new_n584_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1325gat));
  NOR3_X1   g388(.A1(new_n560_), .A2(G15gat), .A3(new_n362_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT100), .Z(new_n591_));
  OAI21_X1  g390(.A(G15gat), .B1(new_n565_), .B2(new_n362_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT41), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(G1326gat));
  INV_X1    g393(.A(new_n372_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G22gat), .B1(new_n565_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT101), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT42), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n598_), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n560_), .A2(G22gat), .A3(new_n595_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(G1327gat));
  NOR2_X1   g401(.A1(new_n558_), .A2(new_n519_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n505_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(G29gat), .B1(new_n605_), .B2(new_n244_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT44), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n559_), .A2(KEYINPUT43), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n559_), .A2(KEYINPUT103), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n610_));
  AOI211_X1 g409(.A(new_n610_), .B(new_n551_), .C1(new_n558_), .C2(new_n550_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n374_), .A2(new_n384_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n564_), .A2(new_n608_), .B1(new_n612_), .B2(KEYINPUT43), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n503_), .A2(new_n518_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT102), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n607_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n564_), .A2(new_n608_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(KEYINPUT43), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n615_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n616_), .A2(new_n621_), .A3(new_n244_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n606_), .B1(new_n622_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g422(.A1(new_n616_), .A2(new_n621_), .A3(new_n569_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G36gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n604_), .A2(G36gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n628_), .B2(new_n569_), .ZN(new_n629_));
  NOR4_X1   g428(.A1(new_n604_), .A2(G36gat), .A3(new_n570_), .A4(new_n626_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n625_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n625_), .A2(new_n631_), .A3(KEYINPUT46), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1329gat));
  NAND4_X1  g435(.A1(new_n616_), .A2(new_n621_), .A3(G43gat), .A4(new_n361_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n604_), .A2(new_n362_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(G43gat), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g439(.A1(new_n616_), .A2(new_n621_), .A3(new_n372_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G50gat), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n595_), .A2(G50gat), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT105), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n605_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n648_), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1331gat));
  INV_X1    g449(.A(new_n502_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n463_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n385_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n519_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n555_), .A2(new_n544_), .A3(new_n557_), .ZN(new_n656_));
  NOR4_X1   g455(.A1(new_n655_), .A2(new_n395_), .A3(new_n561_), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n655_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(KEYINPUT107), .A3(new_n559_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n660_));
  INV_X1    g459(.A(new_n559_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n655_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n659_), .A2(KEYINPUT108), .A3(new_n662_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n244_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n657_), .B1(new_n667_), .B2(new_n395_), .ZN(G1332gat));
  INV_X1    g467(.A(KEYINPUT48), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n655_), .A2(new_n570_), .A3(new_n656_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT109), .B1(new_n670_), .B2(new_n396_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n670_), .A2(KEYINPUT109), .A3(new_n396_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n673_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(KEYINPUT48), .A3(new_n671_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n659_), .A2(new_n396_), .A3(new_n569_), .A4(new_n662_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n676_), .A3(new_n677_), .ZN(G1333gat));
  NAND3_X1  g477(.A1(new_n658_), .A2(new_n361_), .A3(new_n558_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(G71gat), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G71gat), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n362_), .A2(G71gat), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n681_), .A2(new_n682_), .B1(new_n663_), .B2(new_n683_), .ZN(G1334gat));
  NAND3_X1  g483(.A1(new_n658_), .A2(new_n372_), .A3(new_n558_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G78gat), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT50), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT50), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n595_), .A2(G78gat), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n687_), .A2(new_n688_), .B1(new_n663_), .B2(new_n689_), .ZN(G1335gat));
  NAND2_X1  g489(.A1(new_n654_), .A2(new_n603_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n244_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n613_), .A2(new_n519_), .A3(new_n653_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(new_n244_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g495(.A(G92gat), .B1(new_n692_), .B2(new_n569_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n694_), .A2(new_n569_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n429_), .A3(new_n361_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n619_), .A2(new_n518_), .A3(new_n361_), .A4(new_n652_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT111), .B1(new_n701_), .B2(G99gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT51), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(new_n700_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1338gat));
  NAND3_X1  g507(.A1(new_n692_), .A2(new_n409_), .A3(new_n372_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n619_), .A2(new_n518_), .A3(new_n372_), .A4(new_n652_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT52), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G106gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G106gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT53), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT53), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n709_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1339gat));
  NOR2_X1   g517(.A1(new_n569_), .A2(new_n561_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n454_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n452_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n446_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n723_), .A2(new_n725_), .A3(KEYINPUT55), .A4(new_n450_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n453_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n388_), .B1(new_n728_), .B2(new_n445_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n459_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT112), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT56), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n459_), .C1(new_n727_), .C2(new_n729_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n731_), .A2(new_n737_), .A3(new_n732_), .A4(new_n734_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT56), .B(new_n459_), .C1(new_n727_), .C2(new_n729_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n651_), .A3(new_n460_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n487_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n486_), .A2(new_n742_), .A3(new_n489_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n497_), .C1(new_n742_), .C2(new_n492_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n500_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n462_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT114), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n656_), .B1(new_n741_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT57), .B1(new_n749_), .B2(KEYINPUT115), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  INV_X1    g551(.A(new_n739_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n735_), .B2(KEYINPUT113), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n502_), .B1(new_n754_), .B2(new_n738_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n747_), .B1(new_n755_), .B2(new_n460_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n751_), .B(new_n752_), .C1(new_n756_), .C2(new_n656_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n730_), .A2(new_n732_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n460_), .B(new_n745_), .C1(new_n758_), .C2(new_n753_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n661_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n750_), .A2(new_n757_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n518_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n559_), .A2(new_n519_), .A3(new_n502_), .A4(new_n463_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT54), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n720_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n363_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT59), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n766_), .B2(new_n363_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n766_), .A2(KEYINPUT117), .A3(new_n363_), .A4(new_n768_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(G113gat), .A3(new_n651_), .A4(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G113gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n763_), .A2(new_n765_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n363_), .A3(new_n719_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(new_n502_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n775_), .A2(new_n779_), .ZN(G1340gat));
  AOI21_X1  g579(.A(new_n772_), .B1(new_n778_), .B2(KEYINPUT59), .ZN(new_n781_));
  INV_X1    g580(.A(new_n769_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n464_), .B(new_n774_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G120gat), .ZN(new_n784_));
  INV_X1    g583(.A(G120gat), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n785_), .A2(KEYINPUT60), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n463_), .B2(KEYINPUT60), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n766_), .A2(new_n363_), .A3(new_n786_), .A4(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT118), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n784_), .A2(new_n789_), .ZN(G1341gat));
  NAND4_X1  g589(.A1(new_n773_), .A2(G127gat), .A3(new_n519_), .A4(new_n774_), .ZN(new_n791_));
  INV_X1    g590(.A(G127gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n778_), .B2(new_n518_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1342gat));
  NAND4_X1  g593(.A1(new_n773_), .A2(G134gat), .A3(new_n661_), .A4(new_n774_), .ZN(new_n795_));
  INV_X1    g594(.A(G134gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n778_), .B2(new_n558_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1343gat));
  AND3_X1   g597(.A1(new_n766_), .A2(new_n362_), .A3(new_n372_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n651_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n464_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT119), .B(G148gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1345gat));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n519_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT61), .B(G155gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  AOI21_X1  g606(.A(G162gat), .B1(new_n799_), .B2(new_n656_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n609_), .A2(new_n611_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(G162gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n799_), .B2(new_n810_), .ZN(G1347gat));
  NAND2_X1  g610(.A1(new_n569_), .A2(new_n561_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AND4_X1   g612(.A1(new_n651_), .A2(new_n777_), .A3(new_n363_), .A4(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n277_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(KEYINPUT120), .A2(KEYINPUT62), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n814_), .A2(new_n259_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n816_), .B(new_n817_), .C1(new_n814_), .C2(new_n277_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(G1348gat));
  AND2_X1   g622(.A1(new_n777_), .A2(new_n363_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n260_), .A2(KEYINPUT121), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n464_), .A3(new_n813_), .A4(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n260_), .A2(KEYINPUT121), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT122), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n826_), .B(new_n828_), .ZN(G1349gat));
  NAND2_X1  g628(.A1(new_n269_), .A2(KEYINPUT123), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n824_), .A2(new_n813_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n519_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n831_), .A2(new_n519_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n275_), .B1(KEYINPUT123), .B2(new_n274_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(G1350gat));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n273_), .A3(new_n656_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n831_), .A2(new_n661_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n270_), .ZN(G1351gat));
  INV_X1    g637(.A(G197gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT125), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n812_), .A2(new_n361_), .A3(new_n595_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n777_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT124), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n777_), .A2(new_n844_), .A3(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n840_), .B1(new_n846_), .B2(new_n651_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(KEYINPUT125), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n846_), .A2(KEYINPUT125), .A3(new_n839_), .A4(new_n651_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1352gat));
  AND3_X1   g650(.A1(new_n846_), .A2(G204gat), .A3(new_n464_), .ZN(new_n852_));
  AOI21_X1  g651(.A(G204gat), .B1(new_n846_), .B2(new_n464_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1353gat));
  NAND2_X1  g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n846_), .A2(new_n519_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT126), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n858_));
  INV_X1    g657(.A(G211gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n518_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n857_), .A3(new_n858_), .A4(new_n859_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1354gat));
  AOI21_X1  g664(.A(G218gat), .B1(new_n846_), .B2(new_n656_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n559_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(G218gat), .B2(new_n867_), .ZN(G1355gat));
endmodule


