//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_;
  XOR2_X1   g000(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n205_), .A2(KEYINPUT83), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(KEYINPUT83), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n204_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT84), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(KEYINPUT83), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n214_), .A2(KEYINPUT25), .B1(new_n215_), .B2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n217_), .A2(new_n215_), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(new_n219_), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n217_), .B1(new_n215_), .B2(G190gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n209_), .A2(new_n212_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT85), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n209_), .A2(new_n222_), .A3(new_n212_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT23), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n228_), .B1(G183gat), .B2(G190gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n236_), .A2(KEYINPUT86), .A3(G169gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT86), .B1(new_n236_), .B2(G169gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(G176gat), .B1(new_n236_), .B2(G169gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n210_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT30), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(KEYINPUT30), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n202_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n242_), .A2(KEYINPUT30), .ZN(new_n247_));
  INV_X1    g046(.A(new_n202_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT87), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G15gat), .B(G43gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n246_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT90), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n249_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT90), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n246_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT31), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT90), .B(new_n268_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G228gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275_));
  INV_X1    g074(.A(G204gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G197gat), .ZN(new_n277_));
  INV_X1    g076(.A(G197gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G204gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n275_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(G211gat), .A2(G218gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G211gat), .A2(G218gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT94), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT94), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n280_), .A2(new_n286_), .A3(new_n283_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n277_), .A2(new_n279_), .A3(new_n275_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n280_), .A2(new_n283_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n285_), .A2(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT91), .B1(new_n292_), .B2(KEYINPUT1), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(G155gat), .A4(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(KEYINPUT1), .ZN(new_n297_));
  OR2_X1    g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G141gat), .B(G148gat), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI22_X1  g103(.A1(KEYINPUT92), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n304_), .A2(new_n305_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n298_), .A2(new_n292_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n291_), .B1(new_n301_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n274_), .B1(new_n290_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n301_), .A2(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n289_), .A2(new_n288_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n287_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n286_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(new_n320_), .A3(new_n273_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G78gat), .B(G106gat), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(KEYINPUT97), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n301_), .A2(new_n312_), .A3(new_n291_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT28), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n299_), .A2(new_n300_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n291_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G22gat), .B(G50gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(KEYINPUT97), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n314_), .A2(new_n321_), .A3(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n325_), .A2(new_n332_), .A3(new_n334_), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT95), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n322_), .A2(new_n324_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n314_), .A2(new_n321_), .A3(KEYINPUT95), .A4(new_n323_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT96), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(KEYINPUT93), .A3(new_n332_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT93), .ZN(new_n345_));
  INV_X1    g144(.A(new_n332_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(new_n333_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n342_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n343_), .B1(new_n342_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n337_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT98), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT98), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n337_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT25), .B(G183gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n204_), .A2(new_n205_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n233_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n231_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n235_), .A2(new_n210_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n320_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT19), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n241_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n233_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n223_), .B2(KEYINPUT85), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n372_), .B2(new_n226_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n366_), .B(new_n369_), .C1(new_n373_), .C2(new_n290_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT18), .B(G64gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  AND2_X1   g177(.A1(new_n360_), .A2(new_n363_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n379_), .B2(new_n290_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n373_), .B2(new_n290_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n374_), .B(new_n378_), .C1(new_n381_), .C2(new_n369_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT27), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n290_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n368_), .B1(new_n384_), .B2(new_n365_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n234_), .A2(new_n241_), .A3(new_n290_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n364_), .B2(new_n320_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n369_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n378_), .B(KEYINPUT105), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n383_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n378_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n384_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n369_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT27), .B1(new_n396_), .B2(new_n382_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n265_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n266_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n266_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n265_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n315_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n267_), .A2(new_n301_), .A3(new_n312_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n315_), .A2(new_n408_), .A3(new_n404_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n399_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n399_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n410_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n415_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT104), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n398_), .A2(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n272_), .A2(new_n355_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT103), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(KEYINPUT33), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n415_), .C1(new_n410_), .C2(new_n417_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n407_), .A2(new_n399_), .A3(new_n409_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT100), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT100), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n405_), .A2(new_n416_), .A3(new_n406_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n414_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT99), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(KEYINPUT99), .A3(new_n414_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n430_), .A2(new_n431_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n428_), .A2(new_n396_), .A3(new_n382_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT101), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n431_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n430_), .A2(new_n440_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT101), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n382_), .A4(new_n396_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n378_), .A2(KEYINPUT32), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n374_), .B(new_n444_), .C1(new_n381_), .C2(new_n369_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT102), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n390_), .A2(KEYINPUT32), .A3(new_n378_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n395_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(KEYINPUT102), .A3(new_n374_), .A4(new_n444_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n447_), .A2(new_n448_), .A3(new_n420_), .A4(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n439_), .A2(new_n443_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n424_), .B1(new_n452_), .B2(new_n355_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n355_), .A2(new_n421_), .A3(new_n398_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n439_), .A2(new_n443_), .A3(new_n451_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(KEYINPUT103), .A3(new_n352_), .A4(new_n354_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n423_), .B1(new_n457_), .B2(new_n272_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT6), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n460_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT66), .ZN(new_n466_));
  OR2_X1    g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G85gat), .B(G92gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n459_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  AOI211_X1 g272(.A(KEYINPUT8), .B(new_n471_), .C1(new_n469_), .C2(new_n461_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n476_));
  INV_X1    g275(.A(G85gat), .ZN(new_n477_));
  INV_X1    g276(.A(G92gat), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n476_), .A2(KEYINPUT9), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(KEYINPUT9), .B2(new_n476_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT10), .B(G99gat), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n480_), .B(new_n461_), .C1(G106gat), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT67), .B(G71gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G78gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT11), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(KEYINPUT11), .A3(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n483_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n475_), .A2(new_n482_), .A3(new_n490_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n494_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G230gat), .A2(G233gat), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n483_), .A2(KEYINPUT68), .A3(KEYINPUT12), .A4(new_n491_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n495_), .A2(new_n498_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n492_), .A2(new_n496_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G120gat), .B(G148gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G204gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT5), .B(G176gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT70), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n504_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n508_), .B(KEYINPUT69), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT13), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n516_), .A3(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G29gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT15), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  INV_X1    g322(.A(G1gat), .ZN(new_n524_));
  INV_X1    g323(.A(G8gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G8gat), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n521_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT80), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n531_), .B(new_n521_), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(G229gat), .A3(G233gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n518_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n458_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n475_), .A2(new_n482_), .A3(new_n521_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n483_), .A2(new_n522_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n554_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n552_), .B(new_n559_), .C1(new_n554_), .C2(new_n558_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT74), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT36), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT76), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n568_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n562_), .A2(new_n573_), .A3(new_n563_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT75), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n562_), .A2(KEYINPUT75), .A3(new_n563_), .A4(new_n573_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n571_), .A3(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n576_), .A2(new_n577_), .B1(new_n581_), .B2(KEYINPUT37), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n531_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n490_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT16), .B(G183gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n589_), .B(KEYINPUT17), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n585_), .A2(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT79), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT79), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n592_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n582_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n549_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT106), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n421_), .B(KEYINPUT107), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n524_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n576_), .A2(new_n598_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n549_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n421_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n604_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n608_), .A3(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT109), .ZN(new_n611_));
  INV_X1    g410(.A(new_n398_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n549_), .A2(new_n612_), .A3(new_n606_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT108), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n525_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n617_), .B2(KEYINPUT39), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT39), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n615_), .A2(new_n616_), .A3(KEYINPUT109), .A4(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n601_), .A2(new_n525_), .A3(new_n612_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1325gat));
  OAI21_X1  g425(.A(G15gat), .B1(new_n607_), .B2(new_n272_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT41), .Z(new_n628_));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n272_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n601_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(new_n355_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n607_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n601_), .A2(new_n636_), .A3(new_n355_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1327gat));
  NAND2_X1  g437(.A1(new_n576_), .A2(new_n598_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT112), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n549_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT113), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n549_), .A2(KEYINPUT113), .A3(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n421_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n582_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT111), .B1(new_n458_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n458_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n510_), .A2(new_n516_), .A3(new_n513_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n516_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n547_), .B(new_n598_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT110), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(G29gat), .A3(new_n602_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT44), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n648_), .B1(new_n663_), .B2(new_n665_), .ZN(G1328gat));
  NOR2_X1   g465(.A1(new_n398_), .A2(G36gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n646_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT45), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n646_), .A2(new_n670_), .A3(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT114), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n662_), .A2(new_n612_), .A3(new_n665_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(G36gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n612_), .B1(new_n664_), .B2(KEYINPUT44), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n661_), .B(new_n658_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n673_), .B(G36gat), .C1(new_n676_), .C2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n672_), .B1(new_n675_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n672_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  NAND4_X1  g483(.A1(new_n662_), .A2(G43gat), .A3(new_n630_), .A4(new_n665_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n645_), .A2(new_n272_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(G43gat), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g487(.A(G50gat), .B1(new_n646_), .B2(new_n355_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n662_), .A2(G50gat), .A3(new_n355_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n665_), .ZN(G1331gat));
  INV_X1    g490(.A(new_n458_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n518_), .A2(new_n547_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n599_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G57gat), .B1(new_n697_), .B2(new_n602_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n694_), .A2(new_n598_), .A3(new_n576_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n647_), .A2(G57gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(G1332gat));
  INV_X1    g500(.A(G64gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n699_), .B2(new_n612_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n702_), .A3(new_n612_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n699_), .B2(new_n630_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT49), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n709_), .A3(new_n630_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1334gat));
  NAND2_X1  g512(.A1(new_n699_), .A2(new_n355_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G78gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT50), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n633_), .A2(G78gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n696_), .B2(new_n717_), .ZN(G1335gat));
  AND2_X1   g517(.A1(new_n695_), .A2(new_n640_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G85gat), .B1(new_n719_), .B2(new_n602_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n654_), .A2(KEYINPUT116), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n693_), .A2(new_n598_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n654_), .A2(KEYINPUT116), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n421_), .A2(new_n477_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n726_), .B2(new_n727_), .ZN(G1336gat));
  AOI21_X1  g527(.A(G92gat), .B1(new_n719_), .B2(new_n612_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT117), .Z(new_n730_));
  NOR3_X1   g529(.A1(new_n725_), .A2(new_n478_), .A3(new_n398_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n725_), .B2(new_n272_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n272_), .A2(new_n481_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT118), .B1(new_n719_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g536(.A1(new_n654_), .A2(new_n355_), .A3(new_n723_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G106gat), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT52), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(KEYINPUT52), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n633_), .A2(G106gat), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n740_), .A2(new_n741_), .B1(new_n719_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n743_), .B(new_n745_), .ZN(G1339gat));
  NOR2_X1   g545(.A1(new_n655_), .A2(new_n656_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n547_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n599_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n749_), .B(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n501_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n501_), .B2(new_n753_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n495_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n503_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n755_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n512_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n501_), .A2(new_n753_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT55), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n501_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n757_), .A2(new_n503_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n512_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n761_), .A2(new_n547_), .A3(new_n510_), .A4(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n545_), .B1(new_n538_), .B2(new_n536_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n534_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n536_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n546_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n514_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT57), .A3(new_n575_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n761_), .A2(new_n510_), .A3(new_n773_), .A4(new_n768_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT70), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n509_), .B(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n766_), .A2(new_n512_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(KEYINPUT56), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(KEYINPUT58), .A3(new_n773_), .A4(new_n768_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n582_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n776_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT57), .B1(new_n775_), .B2(new_n575_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n598_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n752_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n272_), .A2(new_n355_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n602_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(new_n612_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(KEYINPUT59), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(new_n790_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n790_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n785_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n775_), .A2(new_n575_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n779_), .A2(new_n784_), .A3(KEYINPUT122), .A4(new_n582_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n798_), .A2(new_n801_), .A3(new_n802_), .A4(new_n776_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n598_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n796_), .B1(new_n804_), .B2(new_n752_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n795_), .B(new_n547_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G113gat), .ZN(new_n808_));
  INV_X1    g607(.A(new_n547_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(G113gat), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n805_), .A2(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT123), .B(new_n796_), .C1(new_n804_), .C2(new_n752_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n810_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n808_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT124), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n814_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1340gat));
  OR2_X1    g618(.A1(new_n812_), .A2(new_n813_), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n518_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n820_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n795_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G120gat), .B1(new_n824_), .B2(new_n518_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n824_), .A2(new_n827_), .A3(new_n598_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n820_), .A2(new_n597_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n827_), .ZN(G1342gat));
  INV_X1    g629(.A(G134gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n824_), .A2(new_n831_), .A3(new_n649_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n820_), .A2(new_n576_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n831_), .ZN(G1343gat));
  AOI21_X1  g633(.A(new_n630_), .B1(new_n804_), .B2(new_n752_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n793_), .A2(new_n633_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n809_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n518_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n598_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT61), .B(G155gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  NAND4_X1  g643(.A1(new_n835_), .A2(G162gat), .A3(new_n582_), .A4(new_n836_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n837_), .A2(new_n575_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G162gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT125), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n845_), .B(new_n849_), .C1(new_n846_), .C2(G162gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1347gat));
  NOR2_X1   g650(.A1(new_n602_), .A2(new_n398_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n789_), .A2(new_n790_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT126), .A3(new_n547_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n853_), .B2(new_n809_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(G169gat), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n854_), .A2(new_n547_), .A3(new_n361_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n855_), .A2(KEYINPUT62), .A3(new_n857_), .A4(G169gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(G1348gat));
  AOI21_X1  g662(.A(G176gat), .B1(new_n854_), .B2(new_n747_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n355_), .B1(new_n804_), .B2(new_n752_), .ZN(new_n865_));
  AND4_X1   g664(.A1(G176gat), .A2(new_n747_), .A3(new_n630_), .A4(new_n852_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  NOR3_X1   g666(.A1(new_n853_), .A2(new_n357_), .A3(new_n598_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n865_), .A2(new_n630_), .A3(new_n597_), .A4(new_n852_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n219_), .B2(new_n869_), .ZN(G1350gat));
  OAI21_X1  g669(.A(G190gat), .B1(new_n853_), .B2(new_n649_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n576_), .A2(new_n356_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n853_), .B2(new_n872_), .ZN(G1351gat));
  NOR3_X1   g672(.A1(new_n633_), .A2(new_n647_), .A3(new_n398_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n835_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n809_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n278_), .ZN(G1352gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n518_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1353gat));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n875_), .A2(new_n598_), .A3(new_n881_), .A4(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n875_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n597_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n881_), .ZN(G1354gat));
  AND3_X1   g685(.A1(new_n884_), .A2(G218gat), .A3(new_n582_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G218gat), .B1(new_n884_), .B2(new_n576_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1355gat));
endmodule


