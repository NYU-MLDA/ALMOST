//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT70), .B(G43gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G50gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n205_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n219_));
  AND2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT10), .B(G99gat), .Z(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G85gat), .B(G92gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n229_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n223_), .B(new_n226_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n220_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(KEYINPUT66), .A3(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT7), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n227_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n237_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  AOI211_X1 g049(.A(KEYINPUT8), .B(new_n227_), .C1(new_n223_), .C2(new_n247_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n236_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n215_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n205_), .A2(new_n209_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(new_n236_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n259_), .A2(new_n261_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n254_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(KEYINPUT72), .A3(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n253_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT72), .B1(new_n256_), .B2(new_n262_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT73), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT73), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n271_), .B(new_n264_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n265_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G190gat), .B(G218gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G134gat), .B(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n279_));
  AOI211_X1 g078(.A(new_n279_), .B(new_n265_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n277_), .B(new_n278_), .C1(new_n280_), .C2(new_n276_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n273_), .ZN(new_n283_));
  OAI211_X1 g082(.A(KEYINPUT36), .B(new_n282_), .C1(new_n283_), .C2(new_n279_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT37), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G1gat), .A2(G8gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT76), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT14), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n290_), .B2(KEYINPUT14), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G71gat), .B(G78gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n301_), .B(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n306_), .B2(new_n303_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n300_), .B(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n308_), .A2(KEYINPUT77), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n310_));
  XOR2_X1   g109(.A(G183gat), .B(G211gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(G127gat), .B(G155gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n309_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(KEYINPUT77), .B2(new_n308_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n308_), .B(KEYINPUT79), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n315_), .B(KEYINPUT17), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .A4(KEYINPUT37), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n288_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT80), .ZN(new_n325_));
  INV_X1    g124(.A(new_n307_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n326_), .B(new_n236_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT68), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n252_), .A2(new_n307_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n252_), .A2(KEYINPUT12), .A3(new_n307_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(new_n335_), .A3(new_n328_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(new_n333_), .A3(new_n334_), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n338_), .A3(new_n327_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n328_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n252_), .A2(KEYINPUT67), .A3(new_n307_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT5), .B(G176gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G204gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G120gat), .B(G148gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT13), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n352_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n325_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT81), .ZN(new_n358_));
  INV_X1    g157(.A(G1gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G113gat), .B(G141gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G169gat), .B(G197gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n205_), .A2(new_n209_), .A3(new_n297_), .A4(new_n296_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n215_), .B2(new_n298_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G229gat), .A2(G233gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n210_), .A2(new_n298_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n369_), .A2(new_n364_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n370_), .A2(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n363_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AOI211_X1 g173(.A(KEYINPUT82), .B(new_n362_), .C1(new_n368_), .C2(new_n371_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT83), .Z(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT23), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT86), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n381_), .B2(KEYINPUT24), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT88), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT87), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n381_), .ZN(new_n388_));
  INV_X1    g187(.A(G183gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT25), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT84), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392_));
  INV_X1    g191(.A(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT85), .B(G190gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n392_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n389_), .A2(KEYINPUT25), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n391_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n383_), .A2(new_n388_), .A3(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT89), .B(G176gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G169gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n385_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n379_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n395_), .A2(new_n389_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT30), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(KEYINPUT30), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G127gat), .B(G134gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(new_n412_), .A3(new_n408_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G15gat), .B(G43gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G71gat), .B(G99gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n419_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n415_), .A3(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n420_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n423_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G155gat), .B(G162gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G141gat), .ZN(new_n436_));
  INV_X1    g235(.A(G148gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT91), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT3), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G141gat), .A2(G148gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT2), .Z(new_n441_));
  OAI21_X1  g240(.A(new_n435_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G155gat), .ZN(new_n443_));
  INV_X1    g242(.A(G162gat), .ZN(new_n444_));
  OR3_X1    g243(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT1), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT1), .B1(new_n443_), .B2(new_n444_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n445_), .B(new_n446_), .C1(G155gat), .C2(G162gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n436_), .A2(new_n437_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n440_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT93), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n432_), .B1(new_n452_), .B2(new_n412_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n450_), .B(KEYINPUT93), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n413_), .A2(KEYINPUT101), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n413_), .A2(KEYINPUT101), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n454_), .A2(new_n413_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n431_), .B(new_n453_), .C1(new_n458_), .C2(new_n432_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n431_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G85gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT0), .B(G57gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n460_), .A3(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(KEYINPUT103), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT103), .B1(new_n466_), .B2(new_n468_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT28), .B1(new_n454_), .B2(KEYINPUT29), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n452_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G22gat), .B(G50gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT94), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G211gat), .B(G218gat), .ZN(new_n482_));
  INV_X1    g281(.A(G204gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n483_), .A2(G197gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(G197gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT21), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(KEYINPUT95), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT96), .B1(new_n483_), .B2(G197gat), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n483_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n482_), .B(new_n486_), .C1(new_n490_), .C2(KEYINPUT21), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n482_), .B(KEYINPUT97), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n492_), .A3(KEYINPUT21), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n481_), .B(new_n494_), .C1(new_n452_), .C2(new_n474_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n491_), .A2(new_n493_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n474_), .B1(new_n442_), .B2(new_n449_), .ZN(new_n497_));
  OAI211_X1 g296(.A(G228gat), .B(G233gat), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G78gat), .B(G106gat), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n495_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n472_), .A2(new_n475_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n476_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n477_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n480_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT98), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n477_), .B(new_n505_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT98), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n480_), .A2(new_n502_), .A3(new_n507_), .A4(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n496_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n386_), .B1(G169gat), .B2(G176gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT100), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(KEYINPUT100), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n381_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G190gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(new_n397_), .A3(new_n390_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n380_), .A2(new_n386_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n519_), .A2(new_n379_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n379_), .B1(G183gat), .B2(G190gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n402_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n515_), .B1(new_n494_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n514_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G226gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n406_), .A2(new_n494_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n491_), .A2(new_n493_), .A3(new_n525_), .A4(new_n523_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT20), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n537_), .A3(new_n531_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G8gat), .B(G36gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n232_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT18), .B(G64gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n533_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n528_), .A2(new_n532_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT102), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n536_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n535_), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n534_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n532_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n544_), .B1(new_n550_), .B2(new_n543_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n533_), .A2(new_n538_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n542_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n553_), .A2(new_n544_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT27), .ZN(new_n555_));
  MUX2_X1   g354(.A(new_n551_), .B(new_n554_), .S(new_n555_), .Z(new_n556_));
  AND3_X1   g355(.A1(new_n471_), .A2(new_n513_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT33), .B1(new_n461_), .B2(new_n465_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT33), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n559_), .B(new_n467_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n544_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n458_), .A2(new_n431_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n453_), .B1(new_n458_), .B2(new_n432_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n430_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n467_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n543_), .A2(KEYINPUT32), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n549_), .A2(new_n532_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n545_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n533_), .A2(new_n538_), .A3(new_n567_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n561_), .A2(new_n566_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n513_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n429_), .B1(new_n557_), .B2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n556_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n428_), .A2(new_n471_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n377_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT81), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n325_), .A2(new_n581_), .A3(new_n356_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n358_), .A2(new_n359_), .A3(new_n580_), .A4(new_n582_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n583_), .A2(KEYINPUT104), .A3(new_n471_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT104), .B1(new_n583_), .B2(new_n471_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n575_), .A2(new_n579_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n281_), .A2(new_n284_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT106), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(KEYINPUT106), .A3(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n376_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n355_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT105), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n322_), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G1gat), .B1(new_n599_), .B2(new_n471_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT38), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n588_), .A2(new_n600_), .A3(new_n601_), .ZN(G1324gat));
  NAND3_X1  g401(.A1(new_n358_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n556_), .A2(G8gat), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n556_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n595_), .A2(new_n322_), .A3(new_n607_), .A4(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n608_), .A2(new_n609_), .A3(G8gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n608_), .B2(G8gat), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n606_), .B(KEYINPUT40), .C1(new_n611_), .C2(new_n610_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  OR2_X1    g415(.A1(new_n599_), .A2(new_n429_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(G15gat), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(KEYINPUT41), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(KEYINPUT41), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n603_), .A2(G15gat), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n619_), .B(new_n620_), .C1(new_n429_), .C2(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n599_), .B2(new_n576_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT42), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n576_), .A2(G22gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n603_), .B2(new_n625_), .ZN(G1327gat));
  INV_X1    g425(.A(new_n590_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n321_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n580_), .A2(new_n356_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n471_), .ZN(new_n631_));
  AOI21_X1  g430(.A(G29gat), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n288_), .A2(new_n323_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n589_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT43), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(KEYINPUT44), .A3(new_n321_), .A4(new_n598_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(KEYINPUT43), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n589_), .B2(new_n633_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n321_), .B(new_n598_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n471_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n632_), .B1(new_n644_), .B2(G29gat), .ZN(G1328gat));
  XOR2_X1   g444(.A(new_n556_), .B(KEYINPUT107), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n580_), .A2(new_n356_), .A3(new_n629_), .A4(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(G36gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n636_), .A2(new_n642_), .A3(new_n607_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(G36gat), .ZN(new_n652_));
  OR2_X1    g451(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1329gat));
  XNOR2_X1  g453(.A(KEYINPUT109), .B(G43gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n630_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(new_n429_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n636_), .A2(new_n642_), .A3(G43gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n429_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1330gat));
  NOR3_X1   g460(.A1(new_n643_), .A2(new_n206_), .A3(new_n576_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G50gat), .B1(new_n630_), .B2(new_n513_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1331gat));
  NOR2_X1   g463(.A1(new_n356_), .A2(new_n321_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n595_), .A2(new_n377_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n631_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G57gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n356_), .A2(new_n376_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n589_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n325_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n671_), .A2(G57gat), .A3(new_n471_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1332gat));
  INV_X1    g474(.A(KEYINPUT48), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n666_), .A2(new_n647_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G64gat), .ZN(new_n678_));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT48), .B(new_n679_), .C1(new_n666_), .C2(new_n647_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n647_), .A2(new_n679_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT112), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n678_), .A2(new_n680_), .B1(new_n671_), .B2(new_n682_), .ZN(G1333gat));
  OR3_X1    g482(.A1(new_n671_), .A2(G71gat), .A3(new_n429_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n666_), .A2(new_n428_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT49), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G71gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G71gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1334gat));
  OR3_X1    g488(.A1(new_n671_), .A2(G78gat), .A3(new_n576_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n666_), .A2(new_n513_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(G78gat), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n691_), .B2(G78gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1335gat));
  AND2_X1   g494(.A1(new_n670_), .A2(new_n629_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n631_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n321_), .B(new_n669_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n471_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n699_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g499(.A(G92gat), .B1(new_n696_), .B2(new_n607_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT114), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n698_), .A2(new_n232_), .A3(new_n646_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1337gat));
  OAI21_X1  g503(.A(G99gat), .B1(new_n698_), .B2(new_n429_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(new_n428_), .A3(new_n224_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g507(.A(G106gat), .B1(new_n698_), .B2(new_n576_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n696_), .A2(new_n225_), .A3(new_n513_), .ZN(new_n713_));
  OAI211_X1 g512(.A(G106gat), .B(new_n710_), .C1(new_n698_), .C2(new_n576_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1339gat));
  AND3_X1   g516(.A1(new_n288_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT54), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n356_), .A4(new_n377_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n288_), .A2(new_n322_), .A3(new_n377_), .A4(new_n323_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT54), .B1(new_n721_), .B2(new_n355_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n596_), .A2(new_n349_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n333_), .A2(new_n334_), .A3(new_n327_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n337_), .A2(new_n725_), .B1(new_n726_), .B2(new_n340_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT117), .B1(new_n337_), .B2(new_n725_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n333_), .A2(new_n334_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n327_), .A2(new_n335_), .A3(new_n328_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n335_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n729_), .A2(new_n732_), .A3(new_n733_), .A4(KEYINPUT55), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n727_), .A2(new_n728_), .A3(new_n734_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n735_), .A2(KEYINPUT56), .A3(new_n346_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT56), .B1(new_n735_), .B2(new_n346_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n724_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT118), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n366_), .A2(new_n367_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n370_), .A2(new_n367_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n363_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n372_), .A2(new_n362_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n351_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT118), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n724_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n739_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n590_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n744_), .B(new_n348_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT120), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n735_), .A2(new_n346_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n735_), .A2(KEYINPUT56), .A3(new_n346_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n349_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT120), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(KEYINPUT58), .A4(new_n744_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n752_), .A2(new_n759_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n288_), .A2(new_n323_), .B1(new_n751_), .B2(new_n750_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n749_), .A2(KEYINPUT57), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n748_), .A2(new_n590_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(KEYINPUT119), .A3(new_n764_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n762_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n723_), .B1(new_n769_), .B2(new_n321_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n577_), .A2(new_n429_), .A3(new_n471_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OR3_X1    g571(.A1(new_n770_), .A2(KEYINPUT121), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT121), .B1(new_n770_), .B2(new_n772_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n376_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n748_), .A2(KEYINPUT57), .A3(new_n590_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n750_), .A2(new_n751_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n633_), .A2(new_n778_), .A3(new_n752_), .A4(new_n759_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n321_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n720_), .A2(new_n722_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n772_), .A2(KEYINPUT59), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n780_), .A2(new_n321_), .B1(new_n722_), .B2(new_n720_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n785_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT122), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT59), .B1(new_n770_), .B2(new_n772_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n377_), .ZN(new_n792_));
  AND4_X1   g591(.A1(G113gat), .A2(new_n790_), .A3(new_n791_), .A4(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n776_), .A2(new_n793_), .ZN(G1340gat));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n791_), .A3(new_n355_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT123), .A4(new_n355_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(G120gat), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(G120gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n356_), .B2(KEYINPUT60), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n775_), .B(new_n801_), .C1(KEYINPUT60), .C2(new_n800_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(G1341gat));
  NAND2_X1  g602(.A1(new_n775_), .A2(new_n322_), .ZN(new_n804_));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n790_), .A2(new_n791_), .A3(G127gat), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n804_), .A2(new_n805_), .B1(new_n322_), .B2(new_n806_), .ZN(G1342gat));
  AOI21_X1  g606(.A(G134gat), .B1(new_n775_), .B2(new_n627_), .ZN(new_n808_));
  AND4_X1   g607(.A1(G134gat), .A2(new_n790_), .A3(new_n791_), .A4(new_n633_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n647_), .A2(new_n576_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR4_X1   g611(.A1(new_n770_), .A2(new_n471_), .A3(new_n428_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n376_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n355_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n322_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT61), .B(G155gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1346gat));
  NAND3_X1  g619(.A1(new_n768_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT119), .B1(new_n763_), .B2(new_n764_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n321_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n428_), .B1(new_n823_), .B2(new_n782_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(new_n631_), .A3(new_n633_), .A4(new_n811_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G162gat), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n428_), .B(new_n812_), .C1(new_n823_), .C2(new_n782_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(new_n444_), .A3(new_n631_), .A4(new_n627_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1347gat));
  OR2_X1    g631(.A1(new_n646_), .A2(new_n578_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n787_), .A2(new_n513_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n401_), .A3(new_n376_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n596_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT125), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n576_), .A3(new_n783_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G169gat), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(KEYINPUT62), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT62), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n840_), .B2(new_n841_), .ZN(G1348gat));
  NAND2_X1  g641(.A1(new_n834_), .A2(new_n355_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n770_), .A2(new_n513_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n833_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n845_), .A2(G176gat), .A3(new_n355_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n843_), .A2(new_n400_), .B1(new_n844_), .B2(new_n846_), .ZN(G1349gat));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n322_), .A3(new_n845_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n321_), .B1(new_n397_), .B2(new_n390_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n848_), .A2(new_n389_), .B1(new_n834_), .B2(new_n849_), .ZN(G1350gat));
  NAND3_X1  g649(.A1(new_n834_), .A2(new_n520_), .A3(new_n627_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n834_), .A2(new_n633_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n393_), .ZN(G1351gat));
  NOR2_X1   g652(.A1(new_n631_), .A2(new_n576_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n855_), .B(new_n428_), .C1(new_n823_), .C2(new_n782_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n856_), .A2(new_n647_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n376_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT126), .B(G197gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n376_), .A3(new_n859_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1352gat));
  NAND3_X1  g662(.A1(new_n856_), .A2(new_n355_), .A3(new_n647_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g664(.A1(new_n856_), .A2(new_n322_), .A3(new_n647_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  AND2_X1   g666(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n866_), .B2(new_n867_), .ZN(G1354gat));
  NAND4_X1  g669(.A1(new_n824_), .A2(new_n854_), .A3(new_n633_), .A4(new_n647_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G218gat), .ZN(new_n872_));
  INV_X1    g671(.A(G218gat), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n856_), .A2(new_n873_), .A3(new_n627_), .A4(new_n647_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1355gat));
endmodule


