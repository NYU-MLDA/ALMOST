//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT36), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT10), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT10), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G99gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT64), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT64), .B1(new_n212_), .B2(new_n214_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n210_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(KEYINPUT65), .A3(G85gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n220_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n217_), .A2(new_n219_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G43gat), .B(G50gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G43gat), .B(G50gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n232_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n211_), .A2(new_n210_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT66), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT7), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n227_), .A2(new_n250_), .A3(new_n228_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(KEYINPUT7), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G99gat), .A2(G106gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n246_), .A2(new_n249_), .A3(new_n251_), .A4(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n240_), .B1(new_n255_), .B2(new_n218_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n218_), .A2(new_n240_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n242_), .A2(KEYINPUT66), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n253_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n229_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n257_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n231_), .B(new_n239_), .C1(new_n256_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT73), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(KEYINPUT35), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n231_), .B1(new_n256_), .B2(new_n263_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT15), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n238_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT35), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n271_), .A2(new_n273_), .B1(new_n274_), .B2(new_n268_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n270_), .B1(new_n264_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n264_), .ZN(new_n277_));
  AOI211_X1 g076(.A(new_n274_), .B(new_n268_), .C1(new_n264_), .C2(KEYINPUT73), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n208_), .B(new_n209_), .C1(new_n276_), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n202_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT76), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n209_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n270_), .A2(new_n264_), .A3(new_n275_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n277_), .A2(new_n278_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT75), .B1(new_n288_), .B2(new_n208_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT76), .B1(new_n289_), .B2(new_n202_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n209_), .B(KEYINPUT74), .Z(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n287_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n284_), .A2(new_n290_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G155gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G211gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(KEYINPUT16), .B(G183gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n316_));
  XOR2_X1   g115(.A(G71gat), .B(G78gat), .Z(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n313_), .B(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n302_), .B1(new_n322_), .B2(KEYINPUT17), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(KEYINPUT17), .B2(new_n302_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT77), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n324_), .B(new_n326_), .Z(new_n327_));
  NOR2_X1   g126(.A1(new_n298_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT18), .B(G64gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT20), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT91), .B(G204gat), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G204gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT91), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT91), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G204gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n349_), .B2(G197gat), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n339_), .B(new_n343_), .C1(new_n350_), .C2(new_n340_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G197gat), .A2(G204gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(KEYINPUT21), .B(new_n352_), .C1(new_n341_), .C2(G197gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n343_), .B1(new_n350_), .B2(new_n340_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n354_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT21), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(KEYINPUT93), .A3(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT83), .B(G176gat), .Z(new_n365_));
  INV_X1    g164(.A(G169gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n367_));
  NAND2_X1  g166(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G169gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(KEYINPUT23), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(KEYINPUT23), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G183gat), .A3(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n373_), .B1(new_n377_), .B2(new_n371_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n364_), .B(new_n370_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT25), .B(G183gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G190gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n381_), .A2(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT24), .A3(new_n364_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n386_), .A2(KEYINPUT81), .A3(KEYINPUT24), .A4(new_n364_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n389_), .A3(new_n377_), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n380_), .A2(KEYINPUT85), .A3(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n338_), .B1(new_n363_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n359_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n355_), .A2(KEYINPUT95), .A3(new_n358_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT84), .B1(new_n374_), .B2(new_n376_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n385_), .B(new_n387_), .C1(new_n402_), .C2(new_n373_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n365_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n379_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n377_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n407_), .A3(new_n364_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n401_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n337_), .B1(new_n397_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n394_), .A2(new_n395_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n338_), .B1(new_n359_), .B2(new_n409_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n337_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n334_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G1gat), .B(G29gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G85gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT0), .B(G57gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT99), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT89), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G141gat), .A2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT2), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n430_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(KEYINPUT90), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n426_), .B(new_n427_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G141gat), .B(G148gat), .Z(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n425_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n427_), .B(KEYINPUT1), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G127gat), .A2(G134gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G120gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G127gat), .A2(G134gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(G127gat), .A2(G134gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(G120gat), .B1(new_n449_), .B2(new_n444_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT87), .B(G113gat), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n443_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n437_), .B(new_n442_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(KEYINPUT4), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT98), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT98), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n455_), .A2(new_n461_), .A3(new_n458_), .A4(KEYINPUT4), .ZN(new_n462_));
  AOI211_X1 g261(.A(new_n424_), .B(new_n457_), .C1(new_n460_), .C2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n458_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(new_n423_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n421_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n462_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n457_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n423_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n465_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n421_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n355_), .A2(KEYINPUT93), .A3(new_n358_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT93), .B1(new_n355_), .B2(new_n358_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n396_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n337_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n355_), .A2(new_n358_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(new_n410_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(KEYINPUT20), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n478_), .B2(new_n410_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n474_), .A2(new_n475_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n413_), .B2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n480_), .B(new_n333_), .C1(new_n483_), .C2(new_n337_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n417_), .A2(new_n473_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n472_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n332_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n337_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n476_), .A2(KEYINPUT20), .A3(new_n479_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n480_), .B(new_n332_), .C1(new_n483_), .C2(new_n337_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n469_), .A2(KEYINPUT33), .A3(new_n470_), .A4(new_n471_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n487_), .A2(new_n491_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n464_), .A2(new_n424_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n457_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n471_), .B(new_n495_), .C1(new_n496_), .C2(new_n424_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n485_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499_));
  INV_X1    g298(.A(G227gat), .ZN(new_n500_));
  INV_X1    g299(.A(G233gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n454_), .A2(new_n502_), .ZN(new_n503_));
  OAI22_X1  g302(.A1(new_n452_), .A2(new_n453_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G43gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT31), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G99gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n396_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n394_), .A2(new_n395_), .A3(new_n513_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n509_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n509_), .B1(new_n516_), .B2(new_n515_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n499_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n515_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n516_), .ZN(new_n522_));
  OAI22_X1  g321(.A1(new_n521_), .A2(new_n522_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT88), .A3(new_n517_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n437_), .A2(new_n442_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(G50gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT28), .B(G22gat), .ZN(new_n529_));
  INV_X1    g328(.A(G50gat), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n437_), .A2(new_n442_), .A3(new_n526_), .A4(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n533_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n535_), .B1(new_n539_), .B2(new_n534_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n526_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n399_), .A2(new_n543_), .A3(new_n400_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G228gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n541_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n363_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n540_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n534_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n536_), .A2(new_n538_), .A3(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT96), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(new_n553_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n545_), .A2(new_n547_), .B1(new_n363_), .B2(new_n549_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n552_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n498_), .A2(new_n525_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n523_), .A2(new_n517_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n540_), .A2(new_n551_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n556_), .A2(new_n557_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n552_), .A2(new_n520_), .A3(new_n558_), .A4(new_n524_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n488_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(KEYINPUT27), .A3(new_n492_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT101), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n491_), .A2(new_n492_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT27), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI211_X1 g371(.A(KEYINPUT101), .B(KEYINPUT27), .C1(new_n491_), .C2(new_n492_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n566_), .B(new_n568_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n560_), .B1(new_n574_), .B2(new_n473_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n328_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n249_), .A2(new_n251_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n254_), .B1(new_n583_), .B2(new_n253_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n218_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT8), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n240_), .B(new_n218_), .C1(new_n584_), .C2(new_n229_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n320_), .B1(new_n588_), .B2(new_n231_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT12), .B1(new_n589_), .B2(KEYINPUT68), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n231_), .A3(new_n320_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n271_), .A2(new_n321_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT69), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n600_));
  AOI211_X1 g399(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n271_), .C2(new_n321_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n602_), .A2(KEYINPUT69), .A3(new_n591_), .A4(new_n592_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n581_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n581_), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n605_), .B(new_n608_), .C1(new_n599_), .C2(new_n603_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT71), .ZN(new_n610_));
  OAI22_X1  g409(.A1(new_n607_), .A2(new_n609_), .B1(new_n610_), .B2(KEYINPUT13), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n604_), .A2(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n608_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n604_), .A2(new_n606_), .A3(new_n581_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n239_), .B1(new_n310_), .B2(new_n309_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n311_), .A2(new_n238_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n620_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n238_), .A2(new_n272_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT15), .B1(new_n235_), .B2(new_n237_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n311_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n239_), .A2(new_n310_), .A3(new_n309_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n619_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G169gat), .B(G197gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n632_), .B(KEYINPUT78), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n623_), .B2(new_n628_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT79), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(KEYINPUT79), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT80), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n618_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n576_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n473_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(KEYINPUT102), .A2(KEYINPUT38), .ZN(new_n648_));
  NOR4_X1   g447(.A1(new_n646_), .A2(G1gat), .A3(new_n647_), .A4(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(KEYINPUT102), .A2(KEYINPUT38), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n327_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n575_), .A2(new_n294_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n644_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n618_), .A2(KEYINPUT103), .A3(new_n643_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT104), .Z(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(new_n473_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n651_), .B1(new_n660_), .B2(new_n304_), .ZN(G1324gat));
  OR2_X1    g460(.A1(new_n572_), .A2(new_n573_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n568_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n658_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT39), .ZN(new_n666_));
  INV_X1    g465(.A(new_n646_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n305_), .A3(new_n663_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n525_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n659_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT41), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n559_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n659_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n667_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1327gat));
  AND2_X1   g482(.A1(new_n575_), .A2(new_n296_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n684_), .A2(new_n645_), .A3(new_n327_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n473_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n575_), .A2(new_n687_), .A3(new_n298_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n575_), .A2(new_n298_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n575_), .A2(new_n692_), .A3(new_n687_), .A4(new_n298_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n689_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT106), .B1(new_n657_), .B2(new_n327_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT103), .B1(new_n618_), .B2(new_n643_), .ZN(new_n696_));
  AOI211_X1 g495(.A(new_n654_), .B(new_n642_), .C1(new_n611_), .C2(new_n617_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT106), .B(new_n327_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n694_), .B(KEYINPUT44), .C1(new_n695_), .C2(new_n699_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n473_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n686_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(new_n685_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(G36gat), .A3(new_n664_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n702_), .A2(new_n663_), .A3(new_n703_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G36gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI221_X1 g516(.A(new_n710_), .B1(KEYINPUT110), .B2(KEYINPUT46), .C1(new_n713_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n702_), .A2(G43gat), .A3(new_n561_), .A4(new_n703_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G43gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n707_), .B2(new_n525_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n721_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n722_), .A2(new_n728_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  AOI21_X1  g529(.A(G50gat), .B1(new_n685_), .B2(new_n678_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n559_), .A2(new_n530_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n704_), .B2(new_n732_), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n618_), .A2(new_n643_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n576_), .A2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT112), .Z(new_n736_));
  AOI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n473_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n653_), .A2(new_n734_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n473_), .A2(G57gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(G1332gat));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n741_), .A3(new_n663_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n738_), .B2(new_n663_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n738_), .B2(new_n672_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n736_), .A2(new_n747_), .A3(new_n672_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n738_), .B2(new_n678_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT50), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n736_), .A2(new_n752_), .A3(new_n678_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT114), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n618_), .A2(new_n643_), .A3(new_n652_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n684_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n473_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n694_), .A2(new_n758_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT115), .Z(new_n763_));
  NAND2_X1  g562(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n223_), .B1(new_n647_), .B2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n763_), .B2(new_n765_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n760_), .A2(new_n220_), .A3(new_n663_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n763_), .A2(new_n663_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n220_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n762_), .B2(new_n525_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n561_), .B1(new_n216_), .B2(new_n215_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n759_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n762_), .B2(new_n559_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n694_), .A2(KEYINPUT116), .A3(new_n678_), .A4(new_n758_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(G106gat), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT52), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n775_), .A2(new_n779_), .A3(G106gat), .A4(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n760_), .A2(new_n210_), .A3(new_n678_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(new_n564_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n664_), .A2(new_n473_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT55), .B1(new_n599_), .B2(new_n603_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n590_), .A2(new_n592_), .A3(new_n596_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(G230gat), .A3(G233gat), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n597_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n608_), .B1(new_n792_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT56), .B(new_n608_), .C1(new_n792_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  INV_X1    g601(.A(new_n634_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n619_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n626_), .A2(new_n620_), .A3(new_n627_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n633_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n609_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n614_), .A2(KEYINPUT119), .A3(new_n803_), .A4(new_n806_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT58), .B1(new_n801_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n297_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n296_), .B1(new_n284_), .B2(new_n290_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n791_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n799_), .A2(new_n800_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n298_), .B(KEYINPUT120), .C1(new_n816_), .C2(KEYINPUT58), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n807_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n797_), .A2(KEYINPUT118), .A3(new_n798_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n642_), .A2(new_n609_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n799_), .A2(new_n825_), .A3(new_n800_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n821_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n820_), .B1(new_n827_), .B2(new_n296_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n819_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n821_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n296_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT121), .B1(new_n832_), .B2(KEYINPUT57), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n827_), .A2(new_n834_), .A3(new_n820_), .A4(new_n296_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n652_), .B1(new_n829_), .B2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n328_), .A2(new_n642_), .A3(new_n618_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n328_), .A2(new_n642_), .A3(new_n618_), .A4(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n788_), .B(new_n790_), .C1(new_n837_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n799_), .A2(new_n825_), .A3(new_n800_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n822_), .A2(new_n823_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n831_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT57), .A3(new_n294_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n834_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n294_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n819_), .A3(new_n828_), .A4(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n327_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n843_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n789_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(KEYINPUT122), .A3(new_n788_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n846_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n643_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT59), .B1(new_n856_), .B2(new_n788_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n843_), .B1(new_n853_), .B2(new_n327_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n564_), .A4(new_n789_), .ZN(new_n863_));
  OAI211_X1 g662(.A(G113gat), .B(new_n643_), .C1(new_n860_), .C2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n859_), .A2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g665(.A(new_n446_), .B1(new_n618_), .B2(KEYINPUT60), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n446_), .A2(KEYINPUT60), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n858_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n863_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n844_), .A2(new_n862_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n618_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n446_), .B2(new_n872_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n858_), .B2(new_n652_), .ZN(new_n874_));
  OAI211_X1 g673(.A(G127gat), .B(new_n652_), .C1(new_n860_), .C2(new_n863_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n858_), .B2(new_n296_), .ZN(new_n878_));
  OAI211_X1 g677(.A(G134gat), .B(new_n298_), .C1(new_n860_), .C2(new_n863_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1343gat));
  NOR3_X1   g680(.A1(new_n861_), .A2(new_n565_), .A3(new_n789_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n643_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT123), .B(G141gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1344gat));
  INV_X1    g684(.A(new_n618_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g687(.A1(new_n882_), .A2(new_n652_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  AOI21_X1  g690(.A(G162gat), .B1(new_n882_), .B2(new_n296_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n298_), .A2(G162gat), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT124), .Z(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n882_), .B2(new_n894_), .ZN(G1347gat));
  NOR3_X1   g694(.A1(new_n861_), .A2(new_n473_), .A3(new_n664_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n678_), .A2(new_n525_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n643_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n897_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n643_), .A2(new_n404_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT125), .Z(new_n904_));
  OAI22_X1  g703(.A1(new_n900_), .A2(new_n901_), .B1(new_n902_), .B2(new_n904_), .ZN(G1348gat));
  INV_X1    g704(.A(G176gat), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n902_), .A2(new_n906_), .A3(new_n618_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n902_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n886_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n365_), .B2(new_n909_), .ZN(G1349gat));
  INV_X1    g709(.A(G183gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT126), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n908_), .A2(new_n381_), .A3(new_n652_), .A4(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n902_), .A2(new_n327_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT126), .A2(G183gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n908_), .A2(new_n382_), .A3(new_n296_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G190gat), .B1(new_n902_), .B2(new_n814_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1351gat));
  NOR4_X1   g718(.A1(new_n861_), .A2(new_n473_), .A3(new_n565_), .A4(new_n664_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(G197gat), .A3(new_n643_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n920_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n342_), .B1(new_n924_), .B2(new_n642_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n920_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n643_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n923_), .A2(new_n925_), .A3(new_n926_), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n920_), .A2(new_n886_), .ZN(new_n928_));
  MUX2_X1   g727(.A(new_n349_), .B(G204gat), .S(new_n928_), .Z(G1353gat));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  AND2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n920_), .B(new_n652_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n924_), .A2(new_n327_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n930_), .ZN(G1354gat));
  AOI21_X1  g733(.A(G218gat), .B1(new_n920_), .B2(new_n296_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n298_), .A2(G218gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n920_), .B2(new_n936_), .ZN(G1355gat));
endmodule


