//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n206_), .A2(new_n207_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211_));
  NOR3_X1   g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n211_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G29gat), .B(G36gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT68), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n215_), .B2(new_n208_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT15), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT65), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(KEYINPUT8), .A3(new_n231_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n224_), .A2(new_n225_), .ZN(new_n236_));
  OR2_X1    g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n220_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  INV_X1    g039(.A(G92gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT9), .A3(new_n228_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n236_), .A2(new_n239_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n234_), .A2(new_n235_), .A3(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n211_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n215_), .A2(new_n208_), .A3(new_n213_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n217_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n249_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n235_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT8), .B1(new_n227_), .B2(new_n231_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  AOI211_X1 g056(.A(new_n202_), .B(new_n205_), .C1(new_n251_), .C2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G190gat), .B(G218gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT69), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n205_), .A2(new_n202_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n205_), .A2(new_n202_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n251_), .A2(new_n257_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n269_), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n258_), .B(new_n264_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n262_), .B(KEYINPUT36), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n268_), .B(new_n269_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n258_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n258_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n278_), .B2(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(KEYINPUT37), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT37), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n272_), .A2(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G155gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT16), .ZN(new_n286_));
  XOR2_X1   g085(.A(G183gat), .B(G211gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT17), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  INV_X1    g091(.A(G8gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(G64gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G57gat), .ZN(new_n301_));
  INV_X1    g100(.A(G57gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G64gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT11), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G78gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT66), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT11), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(G71gat), .A2(G78gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G71gat), .A2(G78gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n312_), .B(new_n313_), .C1(new_n314_), .C2(KEYINPUT11), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n306_), .A2(new_n309_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n309_), .B1(new_n306_), .B2(new_n315_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n290_), .B1(new_n299_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n320_), .B2(new_n299_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n289_), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n284_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n317_), .A2(new_n256_), .A3(new_n319_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n316_), .A2(new_n318_), .B1(new_n255_), .B2(new_n254_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G230gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT64), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT12), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n246_), .B(KEYINPUT12), .C1(new_n316_), .C2(new_n318_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n327_), .A4(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G120gat), .B(G148gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(G176gat), .B(G204gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n332_), .A2(new_n337_), .A3(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n348_), .A2(KEYINPUT13), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(KEYINPUT13), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n326_), .A2(KEYINPUT74), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT74), .B1(new_n326_), .B2(new_n351_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT3), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT2), .ZN(new_n361_));
  AOI211_X1 g160(.A(new_n356_), .B(new_n357_), .C1(new_n359_), .C2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n357_), .B1(KEYINPUT1), .B2(new_n355_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(KEYINPUT1), .B2(new_n355_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n358_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n364_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G22gat), .B(G50gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n373_), .B(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G211gat), .B(G218gat), .Z(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G197gat), .B(G204gat), .Z(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n381_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G228gat), .ZN(new_n386_));
  INV_X1    g185(.A(G233gat), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT83), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(KEYINPUT83), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n384_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT85), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n395_), .B(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n376_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n373_), .A2(new_n375_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n373_), .A2(new_n375_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n397_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n401_), .B(new_n402_), .C1(new_n395_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n395_), .A2(new_n403_), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT86), .Z(new_n406_));
  OAI21_X1  g205(.A(new_n400_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT22), .B(G169gat), .ZN(new_n411_));
  INV_X1    g210(.A(G176gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT23), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n413_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT26), .B(G190gat), .Z(new_n422_));
  INV_X1    g221(.A(G183gat), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n423_), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT25), .B1(new_n423_), .B2(KEYINPUT75), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n418_), .A2(new_n414_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n415_), .A2(KEYINPUT23), .ZN(new_n429_));
  INV_X1    g228(.A(G169gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n412_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT24), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .A4(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(KEYINPUT24), .A3(new_n409_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT76), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n421_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT30), .ZN(new_n437_));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT78), .ZN(new_n439_));
  XOR2_X1   g238(.A(G71gat), .B(G99gat), .Z(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n439_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n437_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G127gat), .B(G134gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G113gat), .B(G120gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT31), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n449_), .B(KEYINPUT79), .Z(new_n450_));
  NOR2_X1   g249(.A1(new_n444_), .A2(new_n448_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT80), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n408_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n369_), .A2(KEYINPUT4), .A3(new_n447_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n367_), .A2(KEYINPUT92), .A3(new_n447_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT92), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n367_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n369_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n458_), .B1(new_n461_), .B2(new_n447_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n456_), .B(new_n457_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n462_), .A2(new_n456_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G1gat), .B(G29gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT0), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G57gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT93), .B(G85gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  NAND3_X1  g269(.A1(new_n464_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n471_), .A2(KEYINPUT94), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n419_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n432_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(KEYINPUT89), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT25), .B(G183gat), .Z(new_n477_));
  OAI21_X1  g276(.A(new_n434_), .B1(new_n422_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT88), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(KEYINPUT89), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n428_), .A2(new_n429_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n413_), .B1(new_n482_), .B2(new_n420_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n483_), .A3(new_n385_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT19), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n436_), .B2(new_n384_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n485_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n486_), .A2(new_n489_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT20), .B1(new_n436_), .B2(new_n384_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n481_), .A2(new_n483_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(new_n384_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n496_), .A2(new_n489_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT18), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT91), .ZN(new_n502_));
  XOR2_X1   g301(.A(G64gat), .B(G92gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n455_), .B(new_n457_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n470_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n506_), .B(new_n507_), .C1(new_n455_), .C2(new_n462_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n498_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT94), .B1(new_n471_), .B2(new_n472_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n471_), .A2(new_n472_), .ZN(new_n513_));
  NOR4_X1   g312(.A1(new_n473_), .A2(new_n511_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n464_), .A2(new_n465_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n507_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n516_), .A2(new_n471_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n496_), .A2(new_n489_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT96), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n484_), .A2(new_n491_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n488_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n499_), .A2(KEYINPUT95), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n522_), .A2(KEYINPUT32), .A3(new_n504_), .A4(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n504_), .A2(KEYINPUT32), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n498_), .B2(KEYINPUT95), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n454_), .B1(new_n514_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n505_), .A2(new_n510_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT27), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT98), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT97), .B1(new_n522_), .B2(new_n504_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n519_), .A2(new_n521_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n509_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n536_), .A2(KEYINPUT27), .A3(new_n539_), .A4(new_n505_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n407_), .A2(new_n453_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n407_), .A2(new_n453_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n517_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n528_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n253_), .A2(new_n297_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n297_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n252_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n217_), .A2(new_n551_), .A3(new_n250_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n554_), .B1(new_n557_), .B2(new_n550_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n549_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n549_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n354_), .A2(new_n545_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT99), .ZN(new_n565_));
  INV_X1    g364(.A(new_n517_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n354_), .A2(new_n545_), .A3(new_n567_), .A4(new_n563_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n565_), .A2(new_n292_), .A3(new_n566_), .A4(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n545_), .A2(new_n277_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n351_), .A2(new_n563_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n325_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G1gat), .B1(new_n575_), .B2(new_n517_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(G1324gat));
  INV_X1    g376(.A(KEYINPUT40), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n545_), .A2(new_n277_), .A3(new_n541_), .A4(new_n574_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(G8gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT39), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n582_), .A3(G8gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n565_), .A2(new_n293_), .A3(new_n541_), .A4(new_n568_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT101), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT101), .B1(new_n584_), .B2(new_n585_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n587_), .A2(new_n588_), .A3(KEYINPUT102), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n585_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(new_n586_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n578_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT102), .B1(new_n587_), .B2(new_n588_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n590_), .A3(new_n586_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(KEYINPUT40), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(G1325gat));
  INV_X1    g398(.A(new_n453_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G15gat), .B1(new_n575_), .B2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT41), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT41), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n564_), .A2(G15gat), .A3(new_n600_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(G1326gat));
  OAI21_X1  g404(.A(G22gat), .B1(new_n575_), .B2(new_n407_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT42), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n407_), .A2(G22gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n564_), .B2(new_n608_), .ZN(G1327gat));
  NAND2_X1  g408(.A1(new_n325_), .A2(new_n282_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n573_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n545_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(G29gat), .B1(new_n612_), .B2(new_n566_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n573_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n545_), .A2(new_n284_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n615_), .A2(KEYINPUT43), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(KEYINPUT43), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n614_), .B(new_n325_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n620_), .A2(G29gat), .A3(new_n566_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n619_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n613_), .B1(new_n621_), .B2(new_n622_), .ZN(G1328gat));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n541_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G36gat), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n612_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n541_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n627_), .A2(G36gat), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT45), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT46), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n626_), .A2(KEYINPUT46), .A3(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1329gat));
  NAND4_X1  g434(.A1(new_n620_), .A2(G43gat), .A3(new_n453_), .A4(new_n622_), .ZN(new_n636_));
  INV_X1    g435(.A(G43gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n627_), .B2(new_n600_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n636_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1330gat));
  AOI21_X1  g441(.A(G50gat), .B1(new_n612_), .B2(new_n408_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n620_), .A2(G50gat), .A3(new_n408_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(new_n622_), .ZN(G1331gat));
  NOR2_X1   g444(.A1(new_n351_), .A2(new_n563_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n572_), .A2(new_n324_), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(new_n302_), .A3(new_n517_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT105), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n545_), .A2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n326_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT104), .ZN(new_n652_));
  AOI21_X1  g451(.A(G57gat), .B1(new_n652_), .B2(new_n566_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n649_), .A2(new_n653_), .ZN(G1332gat));
  OAI21_X1  g453(.A(G64gat), .B1(new_n647_), .B2(new_n628_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n541_), .A2(new_n300_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n651_), .B2(new_n658_), .ZN(G1333gat));
  OAI21_X1  g458(.A(G71gat), .B1(new_n647_), .B2(new_n600_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT49), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n600_), .A2(G71gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n651_), .B2(new_n662_), .ZN(G1334gat));
  OAI21_X1  g462(.A(G78gat), .B1(new_n647_), .B2(new_n407_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n407_), .A2(G78gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n651_), .B2(new_n667_), .ZN(G1335gat));
  XNOR2_X1  g467(.A(new_n615_), .B(KEYINPUT43), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n325_), .A3(new_n646_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G85gat), .B1(new_n670_), .B2(new_n517_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n610_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n650_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n240_), .A3(new_n566_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(G1336gat));
  OAI21_X1  g474(.A(G92gat), .B1(new_n670_), .B2(new_n628_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n241_), .A3(new_n541_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1337gat));
  AND2_X1   g477(.A1(new_n237_), .A2(new_n238_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n673_), .A2(new_n679_), .A3(new_n453_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT108), .ZN(new_n681_));
  OAI21_X1  g480(.A(G99gat), .B1(new_n670_), .B2(new_n600_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT51), .ZN(G1338gat));
  XOR2_X1   g483(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n673_), .A2(new_n220_), .A3(new_n408_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n673_), .A2(new_n688_), .A3(new_n220_), .A4(new_n408_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n669_), .A2(new_n408_), .A3(new_n325_), .A4(new_n646_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT52), .B1(new_n691_), .B2(G106gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n685_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n685_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n696_), .A2(new_n692_), .A3(new_n690_), .A4(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n695_), .A2(new_n698_), .ZN(G1339gat));
  NOR2_X1   g498(.A1(new_n541_), .A2(new_n517_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n542_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT112), .Z(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT113), .B(KEYINPUT59), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n280_), .A2(new_n283_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(new_n562_), .A3(new_n351_), .A4(new_n324_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT54), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n346_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n246_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n333_), .B2(new_n328_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n710_), .A2(KEYINPUT55), .A3(new_n335_), .A4(new_n336_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT55), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n337_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n334_), .A2(new_n327_), .A3(new_n336_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n331_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n344_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(KEYINPUT56), .A3(new_n344_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n708_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n557_), .A2(new_n554_), .A3(new_n550_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n550_), .A2(new_n552_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n548_), .B(new_n722_), .C1(new_n723_), .C2(new_n554_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n347_), .A2(new_n559_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n277_), .B1(new_n721_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT111), .ZN(new_n728_));
  INV_X1    g527(.A(new_n346_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n561_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n559_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n716_), .A2(KEYINPUT56), .A3(new_n344_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT56), .B1(new_n716_), .B2(new_n344_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n725_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n277_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT57), .B1(new_n728_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n719_), .A2(new_n720_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n559_), .A2(new_n346_), .A3(new_n724_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT58), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(KEYINPUT58), .A3(new_n740_), .ZN(new_n744_));
  AND4_X1   g543(.A1(new_n283_), .A2(new_n743_), .A3(new_n280_), .A4(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT114), .B1(new_n738_), .B2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n735_), .A2(KEYINPUT57), .A3(new_n277_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n736_), .B1(new_n735_), .B2(new_n277_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT111), .B(new_n282_), .C1(new_n734_), .C2(new_n725_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n284_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n747_), .A3(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n325_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n702_), .B(new_n703_), .C1(new_n707_), .C2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n738_), .A2(new_n745_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n324_), .B1(new_n758_), .B2(new_n747_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n707_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n702_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT59), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n757_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G113gat), .B1(new_n765_), .B2(new_n562_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n562_), .A2(G113gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n762_), .B2(new_n767_), .ZN(G1340gat));
  OAI21_X1  g567(.A(G120gat), .B1(new_n765_), .B2(new_n351_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n351_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT60), .ZN(new_n771_));
  INV_X1    g570(.A(G120gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n763_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n769_), .A2(new_n775_), .ZN(G1341gat));
  OAI21_X1  g575(.A(G127gat), .B1(new_n765_), .B2(new_n325_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n325_), .A2(G127gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n762_), .B2(new_n778_), .ZN(G1342gat));
  INV_X1    g578(.A(G134gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n763_), .A2(new_n780_), .A3(new_n282_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n284_), .B(new_n757_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n783_), .B2(new_n780_), .ZN(G1343gat));
  NOR3_X1   g583(.A1(new_n760_), .A2(new_n453_), .A3(new_n407_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n700_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n562_), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT115), .B(G141gat), .Z(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1344gat));
  INV_X1    g588(.A(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n770_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g591(.A1(new_n786_), .A2(KEYINPUT116), .A3(new_n325_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT116), .B1(new_n786_), .B2(new_n325_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT117), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n797_), .A3(new_n794_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT61), .B(G155gat), .Z(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n796_), .A2(new_n798_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1346gat));
  OAI21_X1  g602(.A(G162gat), .B1(new_n786_), .B2(new_n704_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n277_), .A2(G162gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n786_), .B2(new_n805_), .ZN(G1347gat));
  AOI21_X1  g605(.A(new_n707_), .B1(new_n755_), .B2(new_n325_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n541_), .A2(new_n517_), .A3(new_n453_), .A4(new_n407_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n563_), .A2(new_n411_), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT121), .Z(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n807_), .A2(new_n562_), .A3(new_n808_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n430_), .B1(new_n813_), .B2(KEYINPUT118), .ZN(new_n814_));
  INV_X1    g613(.A(new_n808_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n563_), .C1(new_n756_), .C2(new_n707_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT119), .B(KEYINPUT62), .Z(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n819_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G169gat), .B1(new_n816_), .B2(new_n817_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n813_), .A2(KEYINPUT118), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n822_), .B(new_n824_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n812_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT122), .B(new_n812_), .C1(new_n823_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1348gat));
  AOI21_X1  g632(.A(G176gat), .B1(new_n809_), .B2(new_n770_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n760_), .A2(new_n408_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n628_), .A2(new_n566_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n351_), .A2(new_n412_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n835_), .A2(new_n453_), .A3(new_n836_), .A4(new_n837_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n838_), .A2(KEYINPUT123), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(KEYINPUT123), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n834_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT124), .Z(G1349gat));
  NAND4_X1  g641(.A1(new_n835_), .A2(new_n453_), .A3(new_n324_), .A4(new_n836_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n324_), .A2(new_n477_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n843_), .A2(new_n423_), .B1(new_n809_), .B2(new_n844_), .ZN(G1350gat));
  NAND2_X1  g644(.A1(new_n809_), .A2(new_n284_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G190gat), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT125), .Z(new_n848_));
  NOR4_X1   g647(.A1(new_n807_), .A2(new_n277_), .A3(new_n422_), .A4(new_n808_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1351gat));
  NAND2_X1  g649(.A1(new_n785_), .A2(new_n836_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n563_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G197gat), .ZN(G1352gat));
  XOR2_X1   g653(.A(KEYINPUT126), .B(G204gat), .Z(new_n855_));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G204gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n851_), .A2(new_n351_), .ZN(new_n858_));
  MUX2_X1   g657(.A(new_n855_), .B(new_n857_), .S(new_n858_), .Z(G1353gat));
  NOR2_X1   g658(.A1(new_n851_), .A2(new_n325_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  AND2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n861_), .ZN(G1354gat));
  XOR2_X1   g663(.A(KEYINPUT127), .B(G218gat), .Z(new_n865_));
  NOR3_X1   g664(.A1(new_n851_), .A2(new_n704_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n852_), .A2(new_n282_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1355gat));
endmodule


