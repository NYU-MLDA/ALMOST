//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_;
  AND2_X1   g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n206_), .B(new_n207_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213_));
  AND2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT69), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n203_), .B1(new_n212_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n206_), .A2(new_n207_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT65), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n226_), .B1(new_n233_), .B2(KEYINPUT67), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n206_), .A2(new_n207_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT65), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT65), .B1(new_n230_), .B2(new_n231_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n224_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(G106gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n219_), .B1(new_n248_), .B2(new_n220_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n214_), .B2(KEYINPUT9), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n220_), .A2(KEYINPUT64), .A3(new_n248_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n242_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n255_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n252_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n249_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(KEYINPUT66), .A3(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n241_), .A2(new_n261_), .A3(KEYINPUT70), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n214_), .A2(new_n215_), .A3(new_n213_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT69), .B1(new_n219_), .B2(new_n220_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n225_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n233_), .A2(KEYINPUT67), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n223_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n254_), .A2(new_n260_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n263_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n262_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G57gat), .B(G64gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT11), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT71), .ZN(new_n275_));
  XOR2_X1   g074(.A(G71gat), .B(G78gat), .Z(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(KEYINPUT11), .B2(new_n273_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n272_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n272_), .A2(new_n281_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT72), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(new_n272_), .B2(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n282_), .B1(new_n287_), .B2(KEYINPUT73), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n202_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n283_), .A2(new_n202_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n282_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n241_), .A2(new_n261_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n281_), .A2(new_n295_), .A3(KEYINPUT12), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G120gat), .B(G148gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT5), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G176gat), .B(G204gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n291_), .A2(new_n297_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT13), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n303_), .A2(KEYINPUT13), .A3(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT91), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n319_), .B2(KEYINPUT1), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n316_), .B(new_n320_), .C1(new_n323_), .C2(KEYINPUT1), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n313_), .A2(new_n315_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT93), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329_));
  INV_X1    g128(.A(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT92), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n317_), .A2(new_n334_), .A3(new_n329_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n313_), .A2(new_n315_), .A3(KEYINPUT93), .A4(new_n325_), .ZN(new_n337_));
  OAI22_X1  g136(.A1(new_n317_), .A2(new_n329_), .B1(new_n312_), .B2(new_n325_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n328_), .A2(new_n336_), .A3(new_n337_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT94), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n343_), .A2(KEYINPUT94), .A3(new_n337_), .A4(new_n328_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n323_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n324_), .B1(new_n345_), .B2(KEYINPUT95), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347_));
  AOI211_X1 g146(.A(new_n347_), .B(new_n323_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT29), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G197gat), .B(G204gat), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT21), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G197gat), .B(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT21), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n352_), .A2(new_n355_), .A3(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n349_), .A2(new_n244_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n244_), .B1(new_n349_), .B2(new_n358_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n342_), .A2(new_n344_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n322_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n347_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n345_), .A2(KEYINPUT95), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .A4(new_n324_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G22gat), .B(G50gat), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n371_));
  INV_X1    g170(.A(new_n324_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n364_), .B2(new_n347_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n369_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(new_n366_), .A3(new_n367_), .A4(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n370_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n371_), .B1(new_n370_), .B2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G78gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n376_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n371_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n346_), .A2(new_n348_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n374_), .B1(new_n384_), .B2(new_n366_), .ZN(new_n385_));
  NOR4_X1   g184(.A1(new_n346_), .A2(new_n348_), .A3(KEYINPUT29), .A4(new_n369_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n370_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n382_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n362_), .B1(new_n381_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n380_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n388_), .A3(new_n382_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n361_), .A3(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT25), .B(G183gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT26), .B(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G169gat), .ZN(new_n402_));
  INV_X1    g201(.A(G176gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n404_), .A2(KEYINPUT24), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(KEYINPUT24), .A3(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n396_), .A2(new_n401_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n399_), .A2(new_n409_), .A3(new_n400_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT22), .B(G169gat), .Z(new_n411_));
  OAI211_X1 g210(.A(new_n410_), .B(new_n406_), .C1(new_n411_), .C2(G176gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n358_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT97), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT97), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n358_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT22), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(KEYINPUT87), .B2(new_n402_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n402_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT88), .B(G169gat), .C1(new_n420_), .C2(KEYINPUT87), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n403_), .A3(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n410_), .A2(new_n406_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n407_), .A2(KEYINPUT86), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n396_), .A3(new_n405_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n401_), .B1(KEYINPUT86), .B2(new_n407_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n358_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n419_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n418_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G226gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT19), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G64gat), .B(G92gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT100), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n437_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n358_), .B2(new_n413_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n425_), .A2(new_n426_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n430_), .B2(new_n429_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n358_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n449_), .B2(new_n358_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n445_), .B(new_n447_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n438_), .A2(new_n444_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT104), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT104), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n438_), .A2(new_n457_), .A3(new_n444_), .A4(new_n454_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n418_), .A2(new_n434_), .A3(new_n445_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n453_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n446_), .B1(new_n460_), .B2(new_n451_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n461_), .B2(new_n445_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n444_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT27), .ZN(new_n466_));
  INV_X1    g265(.A(new_n455_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n444_), .B1(new_n438_), .B2(new_n454_), .ZN(new_n468_));
  OR3_X1    g267(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT27), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n390_), .A2(new_n393_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT105), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G134gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G120gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n373_), .A2(new_n367_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(KEYINPUT4), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT101), .Z(new_n482_));
  OAI211_X1 g281(.A(new_n480_), .B(new_n482_), .C1(KEYINPUT4), .C2(new_n479_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G85gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT0), .B(G57gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G15gat), .B(G43gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT89), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT30), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT31), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G227gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(G71gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(G99gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n449_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n496_), .B(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT90), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n476_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n390_), .A2(new_n470_), .A3(new_n393_), .A4(KEYINPUT105), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n473_), .A2(new_n492_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n489_), .A2(KEYINPUT102), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n468_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n455_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n480_), .B(new_n481_), .C1(KEYINPUT4), .C2(new_n479_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n478_), .A2(new_n479_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n488_), .B1(new_n512_), .B2(new_n482_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(KEYINPUT102), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n483_), .A2(new_n484_), .A3(new_n488_), .A4(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n444_), .A2(KEYINPUT32), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT103), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n462_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n462_), .B2(new_n518_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n438_), .A2(new_n454_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n518_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n390_), .A2(new_n393_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT27), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(KEYINPUT27), .B2(new_n465_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n526_), .A2(new_n527_), .B1(new_n530_), .B2(new_n492_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n506_), .B1(new_n531_), .B2(new_n504_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533_));
  INV_X1    g332(.A(G36gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(G29gat), .ZN(new_n535_));
  INV_X1    g334(.A(G29gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(G36gat), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n535_), .A2(new_n537_), .A3(KEYINPUT75), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT75), .B1(new_n535_), .B2(new_n537_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT76), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n536_), .A2(G36gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n534_), .A2(G29gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT76), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n535_), .A2(new_n537_), .A3(KEYINPUT75), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n540_), .A2(new_n541_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n541_), .B1(new_n540_), .B2(new_n548_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n533_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n540_), .A2(new_n548_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n541_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n540_), .A2(new_n548_), .A3(new_n541_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(KEYINPUT15), .A3(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557_));
  INV_X1    g356(.A(G1gat), .ZN(new_n558_));
  INV_X1    g357(.A(G8gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT14), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G8gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n551_), .A2(new_n556_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n554_), .A2(new_n555_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n568_), .A2(KEYINPUT85), .A3(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT85), .B1(new_n568_), .B2(new_n570_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n566_), .B(new_n563_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n570_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n575_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n311_), .A2(new_n532_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT81), .B(KEYINPUT36), .Z(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n262_), .A2(new_n271_), .A3(new_n566_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT34), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n262_), .A2(new_n271_), .A3(KEYINPUT79), .A4(new_n566_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n551_), .B(new_n556_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT77), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT77), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n295_), .A2(new_n599_), .A3(new_n556_), .A4(new_n551_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n592_), .A2(new_n593_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n586_), .B1(new_n596_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT80), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n587_), .A2(new_n588_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n595_), .A2(new_n594_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n598_), .A2(new_n600_), .A3(KEYINPUT78), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT78), .B1(new_n598_), .B2(new_n600_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n589_), .A2(KEYINPUT80), .A3(new_n594_), .A4(new_n595_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n605_), .B1(new_n614_), .B2(new_n602_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT82), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n596_), .A2(new_n604_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n614_), .B2(new_n602_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n584_), .B(KEYINPUT36), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(KEYINPUT83), .A2(KEYINPUT37), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT83), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n617_), .A2(new_n622_), .A3(new_n623_), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n614_), .A2(new_n602_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n605_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n616_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT82), .B(new_n605_), .C1(new_n614_), .C2(new_n602_), .ZN(new_n631_));
  OAI22_X1  g430(.A1(new_n630_), .A2(new_n631_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT16), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n280_), .B(new_n564_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n641_), .B2(KEYINPUT84), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT17), .B1(new_n641_), .B2(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT17), .B(new_n638_), .C1(new_n641_), .C2(KEYINPUT84), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n634_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n581_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n492_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n558_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n532_), .A2(new_n632_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n310_), .A2(new_n647_), .A3(new_n579_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n492_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n652_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n653_), .A2(new_n657_), .A3(new_n658_), .ZN(G1324gat));
  NAND3_X1  g458(.A1(new_n649_), .A2(new_n559_), .A3(new_n529_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G8gat), .B1(new_n656_), .B2(new_n470_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g464(.A(new_n504_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G15gat), .B1(new_n656_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT41), .Z(new_n668_));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n649_), .A2(new_n669_), .A3(new_n504_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1326gat));
  XOR2_X1   g470(.A(new_n527_), .B(KEYINPUT106), .Z(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G22gat), .B1(new_n656_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT42), .ZN(new_n675_));
  INV_X1    g474(.A(G22gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n649_), .A2(new_n676_), .A3(new_n672_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1327gat));
  NOR3_X1   g477(.A1(new_n310_), .A2(new_n646_), .A3(new_n579_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n532_), .A2(new_n680_), .A3(new_n634_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n532_), .B2(new_n634_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n679_), .B(KEYINPUT44), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n492_), .A2(new_n536_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n632_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n647_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n581_), .A2(new_n650_), .A3(new_n691_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n687_), .A2(new_n688_), .B1(new_n536_), .B2(new_n692_), .ZN(G1328gat));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n685_), .A2(new_n529_), .A3(new_n686_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n581_), .A2(new_n534_), .A3(new_n529_), .A4(new_n691_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT45), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n694_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n695_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT107), .B1(new_n695_), .B2(G36gat), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n702_), .B(new_n694_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n703_), .A2(new_n707_), .ZN(G1329gat));
  NAND3_X1  g507(.A1(new_n687_), .A2(G43gat), .A3(new_n504_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n581_), .A2(new_n691_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(new_n666_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(G43gat), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g512(.A(new_n527_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n687_), .A2(G50gat), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n710_), .B2(new_n673_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1331gat));
  NOR3_X1   g517(.A1(new_n311_), .A2(new_n647_), .A3(new_n580_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n654_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n492_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n532_), .A2(new_n579_), .A3(new_n310_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n648_), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n650_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n721_), .A2(new_n725_), .ZN(G1332gat));
  INV_X1    g525(.A(G64gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n727_), .A3(new_n529_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n720_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n529_), .ZN(new_n730_));
  XOR2_X1   g529(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(G64gat), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n723_), .A2(new_n498_), .A3(new_n504_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n729_), .A2(new_n504_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(G71gat), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G71gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1334gat));
  OAI21_X1  g541(.A(G78gat), .B1(new_n720_), .B2(new_n673_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT50), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n723_), .A2(new_n379_), .A3(new_n672_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  NAND3_X1  g545(.A1(new_n310_), .A2(new_n647_), .A3(new_n579_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n492_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n722_), .A2(new_n691_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n217_), .A3(new_n650_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n749_), .B2(new_n470_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n218_), .A3(new_n529_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1337gat));
  NAND4_X1  g555(.A1(new_n751_), .A2(new_n243_), .A3(new_n245_), .A4(new_n504_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G99gat), .B1(new_n749_), .B2(new_n666_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT112), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n759_), .B(new_n761_), .ZN(G1338gat));
  OAI21_X1  g561(.A(KEYINPUT113), .B1(new_n749_), .B2(new_n527_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n532_), .A2(new_n634_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT43), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n532_), .A2(new_n634_), .A3(new_n680_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n747_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n714_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n763_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT52), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n763_), .A2(new_n769_), .A3(new_n772_), .A4(G106gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n751_), .A2(new_n244_), .A3(new_n714_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n774_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1339gat));
  INV_X1    g580(.A(G113gat), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n310_), .A2(new_n580_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n648_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT54), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n648_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n294_), .A2(new_n296_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n202_), .B1(new_n287_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n297_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n292_), .A2(KEYINPUT55), .A3(new_n294_), .A4(new_n296_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n302_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n796_), .B(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n305_), .A2(new_n580_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .A4(new_n578_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n578_), .B1(new_n573_), .B2(new_n569_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n799_), .A2(new_n800_), .B1(new_n306_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n632_), .B1(KEYINPUT116), .B2(KEYINPUT57), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n789_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n306_), .A2(new_n804_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n796_), .B1(new_n797_), .B2(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n795_), .A2(new_n302_), .A3(new_n798_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n580_), .A3(new_n305_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n632_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n795_), .A2(new_n816_), .A3(new_n302_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n815_), .A2(new_n305_), .A3(new_n804_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n819_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n634_), .A3(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n647_), .B1(new_n814_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n788_), .A2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n473_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n650_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n492_), .B1(new_n788_), .B2(new_n823_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT117), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(new_n580_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n825_), .A3(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n826_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n580_), .A2(G113gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT119), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n782_), .A2(new_n832_), .B1(new_n838_), .B2(new_n840_), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n837_), .B2(new_n311_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n828_), .A2(new_n831_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT60), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n310_), .A2(new_n844_), .ZN(new_n845_));
  MUX2_X1   g644(.A(new_n845_), .B(new_n844_), .S(G120gat), .Z(new_n846_));
  OAI21_X1  g645(.A(new_n842_), .B1(new_n843_), .B2(new_n846_), .ZN(G1341gat));
  OAI21_X1  g646(.A(G127gat), .B1(new_n837_), .B2(new_n647_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n647_), .A2(G127gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n843_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n828_), .A2(new_n689_), .A3(new_n831_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n634_), .A2(G134gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT120), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n851_), .A2(new_n852_), .B1(new_n838_), .B2(new_n854_), .ZN(G1343gat));
  NOR3_X1   g654(.A1(new_n527_), .A2(new_n504_), .A3(new_n529_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n829_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n580_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n310_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT121), .B(G148gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1345gat));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n646_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  NAND3_X1  g664(.A1(new_n829_), .A2(new_n689_), .A3(new_n856_), .ZN(new_n866_));
  INV_X1    g665(.A(G162gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n868_), .A2(KEYINPUT122), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(KEYINPUT122), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n627_), .B2(new_n633_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n870_), .B1(new_n857_), .B2(new_n871_), .ZN(G1347gat));
  NOR3_X1   g671(.A1(new_n666_), .A2(new_n650_), .A3(new_n470_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n788_), .B2(new_n823_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n875_), .A2(new_n673_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n411_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n580_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n873_), .A2(new_n580_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT123), .Z(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n672_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n402_), .B1(new_n824_), .B2(new_n881_), .ZN(new_n882_));
  OR2_X1    g681(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n883_));
  NAND2_X1  g682(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n878_), .B(new_n885_), .C1(new_n883_), .C2(new_n882_), .ZN(G1348gat));
  NAND3_X1  g685(.A1(new_n875_), .A2(new_n310_), .A3(new_n673_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n403_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(KEYINPUT125), .A3(new_n403_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n873_), .A2(G176gat), .A3(new_n527_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n311_), .A2(new_n892_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n890_), .A2(new_n891_), .B1(new_n824_), .B2(new_n893_), .ZN(G1349gat));
  NOR2_X1   g693(.A1(new_n647_), .A2(new_n394_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n875_), .A2(new_n673_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n714_), .A2(new_n647_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n824_), .A2(new_n897_), .A3(new_n873_), .A4(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(G183gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n897_), .B1(new_n875_), .B2(new_n898_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n896_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT127), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n896_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1350gat));
  NAND2_X1  g706(.A1(new_n876_), .A2(new_n634_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G190gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n876_), .A2(new_n689_), .A3(new_n395_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1351gat));
  NAND4_X1  g710(.A1(new_n714_), .A2(new_n666_), .A3(new_n492_), .A4(new_n529_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n788_), .B2(new_n823_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n580_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n310_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n646_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n913_), .A2(new_n923_), .A3(new_n689_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n913_), .A2(new_n634_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1355gat));
endmodule


