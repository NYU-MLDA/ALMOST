//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n211_), .C1(KEYINPUT9), .C2(new_n210_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT67), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n214_), .A3(KEYINPUT65), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT7), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT7), .B1(new_n220_), .B2(new_n221_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n214_), .A3(KEYINPUT64), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n209_), .A2(KEYINPUT66), .A3(new_n210_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  INV_X1    g027(.A(new_n210_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(new_n208_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n218_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n234_), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n235_), .B2(KEYINPUT64), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT7), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n236_), .A2(new_n207_), .A3(new_n224_), .A4(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n231_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n218_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n216_), .B1(new_n232_), .B2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(G57gat), .A2(G64gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G57gat), .A2(G64gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n246_));
  INV_X1    g045(.A(G71gat), .ZN(new_n247_));
  INV_X1    g046(.A(G78gat), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n245_), .A2(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G71gat), .A2(G78gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT11), .B1(new_n243_), .B2(new_n244_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT68), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(KEYINPUT11), .C1(new_n243_), .C2(new_n244_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n249_), .A2(new_n250_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n248_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G57gat), .B(G64gat), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n250_), .B(new_n256_), .C1(new_n257_), .C2(KEYINPUT11), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n257_), .B2(KEYINPUT11), .ZN(new_n259_));
  INV_X1    g058(.A(new_n254_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n202_), .B1(new_n242_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT72), .ZN(new_n264_));
  INV_X1    g063(.A(new_n216_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n240_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n255_), .A2(new_n261_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n202_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n264_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n262_), .A2(KEYINPUT70), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n202_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT71), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n268_), .A2(new_n274_), .A3(new_n276_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G230gat), .A2(G233gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n242_), .A2(new_n262_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n273_), .A2(new_n281_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n270_), .A2(new_n283_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n282_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT69), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G120gat), .B(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(G204gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT5), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(KEYINPUT69), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n284_), .A2(new_n288_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n284_), .A2(new_n288_), .A3(new_n295_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n294_), .B(KEYINPUT73), .Z(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT13), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G229gat), .A2(G233gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G1gat), .A2(G8gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT14), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G15gat), .A2(G22gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(G15gat), .A2(G22gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT77), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(KEYINPUT77), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G8gat), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G29gat), .B(G36gat), .Z(new_n316_));
  INV_X1    g115(.A(G43gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G29gat), .B(G36gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G43gat), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(G50gat), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(G50gat), .B1(new_n318_), .B2(new_n320_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n315_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n315_), .A2(new_n323_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n302_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT15), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n318_), .A2(new_n320_), .ZN(new_n330_));
  INV_X1    g129(.A(G50gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n318_), .A2(G50gat), .A3(new_n320_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT15), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n324_), .B(new_n301_), .C1(new_n336_), .C2(new_n315_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n327_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G141gat), .ZN(new_n339_));
  INV_X1    g138(.A(G169gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(KEYINPUT80), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n338_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n300_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT25), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT25), .B(G183gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n348_), .B(new_n351_), .C1(new_n352_), .C2(new_n349_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n340_), .A2(new_n293_), .A3(KEYINPUT82), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(G169gat), .B2(G176gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n340_), .A2(new_n293_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(KEYINPUT24), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364_));
  NAND3_X1  g163(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(KEYINPUT23), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n354_), .A2(new_n356_), .A3(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n353_), .A2(new_n360_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G169gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n358_), .B1(new_n372_), .B2(new_n293_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n363_), .A2(KEYINPUT23), .A3(new_n365_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n361_), .A2(new_n364_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(new_n247_), .ZN(new_n382_));
  INV_X1    g181(.A(G113gat), .ZN(new_n383_));
  OR2_X1    g182(.A1(G127gat), .A2(G134gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G127gat), .A2(G134gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(G120gat), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G120gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n386_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n382_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n381_), .B(G71gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n389_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G43gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G99gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n400_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n393_), .A2(new_n396_), .A3(new_n403_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G141gat), .B(G148gat), .Z(new_n410_));
  NOR2_X1   g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT85), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT1), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n410_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n411_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT2), .ZN(new_n418_));
  INV_X1    g217(.A(G141gat), .ZN(new_n419_));
  INV_X1    g218(.A(G148gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n426_), .A3(new_n413_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n415_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n395_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n415_), .A2(new_n389_), .A3(new_n392_), .A4(new_n427_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n409_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(KEYINPUT4), .A3(new_n430_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n429_), .A2(KEYINPUT93), .A3(KEYINPUT4), .A4(new_n430_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n429_), .A2(KEYINPUT4), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n431_), .B1(new_n438_), .B2(new_n409_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G1gat), .B(G29gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(new_n433_), .B2(new_n432_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n408_), .B1(new_n447_), .B2(new_n435_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n448_), .B2(new_n431_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n407_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n453_), .A2(G36gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(G64gat), .B(G92gat), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(G36gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n456_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT92), .B(G8gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n453_), .B(G36gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n455_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n465_), .B2(new_n458_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT19), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G197gat), .B(G204gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT21), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT21), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(KEYINPUT88), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n472_), .B(KEYINPUT89), .C1(new_n474_), .C2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G211gat), .B(G218gat), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G197gat), .B(G204gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT21), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n486_), .A2(new_n482_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n483_), .B1(new_n487_), .B2(new_n478_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n367_), .ZN(new_n489_));
  AND3_X1   g288(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n492_), .B2(new_n364_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n373_), .B1(new_n493_), .B2(new_n377_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n375_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n492_), .B2(KEYINPUT23), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n348_), .A2(new_n352_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n369_), .A2(new_n340_), .A3(new_n293_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n496_), .A2(new_n360_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n471_), .B1(new_n488_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n478_), .B1(new_n486_), .B2(new_n482_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n477_), .A2(new_n479_), .B1(KEYINPUT21), .B2(new_n481_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n379_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n470_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(new_n499_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n378_), .B(new_n371_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n509_));
  AND4_X1   g308(.A1(KEYINPUT20), .A2(new_n508_), .A3(new_n470_), .A4(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n468_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n462_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n465_), .A2(new_n461_), .A3(new_n458_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n512_), .A2(KEYINPUT97), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT97), .B1(new_n512_), .B2(new_n513_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n470_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n518_));
  AND4_X1   g317(.A1(KEYINPUT20), .A2(new_n508_), .A3(new_n517_), .A4(new_n509_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n511_), .A2(new_n520_), .A3(KEYINPUT27), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n494_), .B(new_n499_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n505_), .A2(KEYINPUT20), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n517_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n371_), .A2(new_n378_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n471_), .B1(new_n488_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n470_), .A3(new_n508_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n527_), .A3(new_n467_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT27), .B1(new_n511_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT98), .B1(new_n521_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT27), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n524_), .A2(new_n527_), .A3(new_n467_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n467_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n511_), .A2(new_n520_), .A3(KEYINPUT27), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT98), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n428_), .A2(KEYINPUT29), .ZN(new_n539_));
  XOR2_X1   g338(.A(G22gat), .B(G50gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT28), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n539_), .B(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G78gat), .B(G106gat), .Z(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(KEYINPUT90), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n543_), .B2(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n428_), .A2(KEYINPUT29), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n504_), .A2(new_n546_), .A3(KEYINPUT87), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G228gat), .A2(G233gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT86), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n547_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n550_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n552_), .B(new_n544_), .C1(new_n543_), .C2(new_n542_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n452_), .B1(new_n538_), .B2(new_n555_), .ZN(new_n556_));
  AOI211_X1 g355(.A(KEYINPUT99), .B(new_n554_), .C1(new_n530_), .C2(new_n537_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n451_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n446_), .B(new_n559_), .C1(new_n448_), .C2(new_n431_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n434_), .A2(new_n437_), .A3(new_n408_), .A4(new_n435_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n429_), .A2(new_n409_), .A3(new_n430_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n565_), .A2(new_n444_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n511_), .A2(new_n567_), .A3(new_n528_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT96), .B1(new_n563_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n468_), .A2(KEYINPUT32), .ZN(new_n572_));
  INV_X1    g371(.A(new_n518_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n519_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n554_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n563_), .A2(KEYINPUT96), .A3(new_n569_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n571_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n534_), .A2(new_n535_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n554_), .B1(new_n581_), .B2(new_n450_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n407_), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n347_), .B1(new_n558_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n268_), .A2(new_n335_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n242_), .A2(new_n323_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n588_), .A2(KEYINPUT35), .A3(new_n590_), .A4(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT35), .A3(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n587_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n590_), .A2(KEYINPUT35), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G134gat), .ZN(new_n600_));
  INV_X1    g399(.A(G162gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(KEYINPUT36), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT75), .Z(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(new_n596_), .A3(new_n593_), .A4(new_n595_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(KEYINPUT37), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n597_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n593_), .A2(new_n595_), .A3(KEYINPUT76), .A4(new_n596_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n603_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n607_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT79), .B(G127gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT70), .A3(KEYINPUT17), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(KEYINPUT17), .B2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n269_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n315_), .ZN(new_n625_));
  MUX2_X1   g424(.A(new_n621_), .B(new_n622_), .S(new_n625_), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n584_), .A2(new_n614_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n450_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n627_), .A2(G1gat), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n629_), .A2(KEYINPUT100), .A3(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n300_), .A2(new_n346_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n558_), .A2(new_n583_), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n612_), .A2(new_n632_), .A3(new_n626_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n450_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n629_), .A2(new_n630_), .B1(G1gat), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT100), .B1(new_n629_), .B2(new_n630_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n631_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT101), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n631_), .A2(new_n640_), .A3(new_n636_), .A4(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1324gat));
  OR3_X1    g441(.A1(new_n627_), .A2(G8gat), .A3(new_n538_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n538_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n634_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G8gat), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1325gat));
  AND2_X1   g450(.A1(new_n405_), .A2(new_n406_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n634_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G15gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  NOR3_X1   g454(.A1(new_n627_), .A2(G15gat), .A3(new_n407_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT102), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n634_), .A2(new_n554_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G22gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT103), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n627_), .A2(G22gat), .A3(new_n555_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n612_), .A2(new_n626_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n584_), .A2(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n668_), .A2(G29gat), .A3(new_n628_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n607_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n612_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(KEYINPUT37), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n652_), .A2(new_n628_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n534_), .A2(new_n536_), .A3(new_n535_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n536_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n555_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT99), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n538_), .A2(new_n452_), .A3(new_n555_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n673_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n582_), .A2(new_n407_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT96), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n681_), .B(new_n568_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n570_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n683_), .B2(new_n578_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n672_), .B1(new_n679_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n626_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT104), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n672_), .B(new_n690_), .C1(new_n679_), .C2(new_n684_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n687_), .A2(new_n688_), .A3(new_n632_), .A4(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(KEYINPUT44), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n614_), .B1(new_n558_), .B2(new_n583_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n686_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n691_), .B(new_n688_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n693_), .A2(KEYINPUT44), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n693_), .A2(KEYINPUT44), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n697_), .A2(new_n347_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n450_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n669_), .B1(new_n701_), .B2(G29gat), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT106), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n538_), .B(KEYINPUT107), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n584_), .A2(new_n704_), .A3(new_n667_), .A4(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT45), .Z(new_n708_));
  OAI21_X1  g507(.A(new_n644_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G36gat), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n710_), .B(new_n712_), .ZN(G1329gat));
  NOR2_X1   g512(.A1(new_n407_), .A2(new_n317_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT109), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n714_), .C1(new_n694_), .C2(new_n700_), .ZN(new_n718_));
  XOR2_X1   g517(.A(KEYINPUT110), .B(G43gat), .Z(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n668_), .B2(new_n407_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n718_), .A3(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT112), .Z(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n716_), .A2(new_n723_), .A3(new_n718_), .A4(new_n720_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1330gat));
  OAI21_X1  g526(.A(new_n554_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n728_), .A2(KEYINPUT113), .A3(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT113), .B1(new_n728_), .B2(G50gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n554_), .A2(new_n331_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT114), .Z(new_n732_));
  OAI22_X1  g531(.A1(new_n729_), .A2(new_n730_), .B1(new_n668_), .B2(new_n732_), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n300_), .A2(new_n346_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n633_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n614_), .A3(new_n626_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n450_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739_));
  OAI21_X1  g538(.A(G57gat), .B1(new_n628_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n612_), .A3(new_n626_), .ZN(new_n741_));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(KEYINPUT115), .B2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n738_), .B1(new_n740_), .B2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n741_), .B2(new_n705_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT116), .B(KEYINPUT117), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT48), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n745_), .B(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n736_), .A2(G64gat), .A3(new_n705_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1333gat));
  NAND3_X1  g549(.A1(new_n737_), .A2(new_n247_), .A3(new_n652_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G71gat), .B1(new_n741_), .B2(new_n407_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT49), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT49), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n741_), .B2(new_n555_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n737_), .A2(new_n248_), .A3(new_n554_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1335gat));
  INV_X1    g558(.A(new_n697_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n734_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n450_), .A2(G85gat), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT118), .Z(new_n763_));
  NAND2_X1  g562(.A1(new_n735_), .A2(new_n667_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n628_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n761_), .A2(new_n763_), .B1(new_n765_), .B2(G85gat), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT119), .Z(G1336gat));
  INV_X1    g566(.A(new_n764_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G92gat), .B1(new_n768_), .B2(new_n644_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n761_), .A2(new_n705_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n761_), .B2(new_n407_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n213_), .A3(new_n652_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n772_), .B(new_n773_), .C1(KEYINPUT120), .C2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT120), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n214_), .A3(new_n554_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n554_), .A3(new_n734_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g584(.A(new_n346_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n300_), .A2(new_n614_), .A3(new_n626_), .A4(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n296_), .A2(new_n346_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n296_), .A2(new_n346_), .A3(KEYINPUT121), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n298_), .ZN(new_n795_));
  AND4_X1   g594(.A1(new_n282_), .A2(new_n273_), .A3(new_n283_), .A4(new_n281_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n271_), .B1(new_n270_), .B2(new_n202_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT72), .B(KEYINPUT12), .C1(new_n268_), .C2(new_n269_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n283_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n281_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n286_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n796_), .B1(KEYINPUT55), .B2(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n264_), .A2(new_n272_), .B1(new_n242_), .B2(new_n262_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n803_), .A2(KEYINPUT55), .A3(new_n282_), .A4(new_n281_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n795_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n282_), .B1(new_n803_), .B2(new_n281_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n284_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n804_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n794_), .B1(new_n808_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n301_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n324_), .B(new_n302_), .C1(new_n336_), .C2(new_n315_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n343_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT122), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n327_), .A2(new_n337_), .A3(new_n344_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT122), .A4(new_n343_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n299_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n612_), .B1(new_n814_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT57), .B(new_n612_), .C1(new_n814_), .C2(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n296_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n822_), .A2(KEYINPUT123), .A3(new_n296_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n795_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n807_), .B(new_n298_), .C1(new_n811_), .C2(new_n804_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n832_), .B(KEYINPUT58), .C1(new_n833_), .C2(new_n834_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n672_), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n827_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n789_), .B1(new_n840_), .B2(new_n688_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n628_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n841_), .A2(new_n407_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n346_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n688_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n789_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n407_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n842_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n841_), .A2(new_n850_), .A3(new_n407_), .A4(new_n843_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n786_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n845_), .B1(new_n854_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g654(.A(new_n390_), .B1(new_n300_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n844_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n390_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n300_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n390_), .ZN(G1341gat));
  AOI21_X1  g658(.A(KEYINPUT59), .B1(new_n848_), .B2(new_n842_), .ZN(new_n860_));
  OAI211_X1 g659(.A(G127gat), .B(new_n626_), .C1(new_n860_), .C2(new_n852_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n862_), .B(new_n863_), .C1(new_n849_), .C2(new_n688_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n841_), .A2(new_n688_), .A3(new_n407_), .A4(new_n843_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT124), .B1(new_n865_), .B2(G127gat), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n861_), .A2(new_n864_), .A3(new_n866_), .ZN(G1342gat));
  AOI21_X1  g666(.A(G134gat), .B1(new_n844_), .B2(new_n671_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n614_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n652_), .A2(new_n555_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n841_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n706_), .A2(new_n628_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n786_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n419_), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n300_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n420_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n688_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  NOR3_X1   g681(.A1(new_n875_), .A2(new_n601_), .A3(new_n614_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n873_), .A2(new_n671_), .A3(new_n874_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n601_), .B2(new_n884_), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n705_), .A2(new_n450_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n848_), .A2(new_n555_), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887_), .B2(new_n786_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n786_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n372_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT62), .B(G169gat), .C1(new_n887_), .C2(new_n786_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  OR3_X1    g693(.A1(new_n887_), .A2(new_n293_), .A3(new_n300_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n293_), .B1(new_n887_), .B2(new_n300_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1349gat));
  NOR3_X1   g696(.A1(new_n887_), .A2(new_n688_), .A3(new_n352_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n887_), .A2(new_n688_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n350_), .B2(new_n899_), .ZN(G1350gat));
  INV_X1    g699(.A(new_n348_), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n887_), .A2(new_n612_), .A3(new_n901_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n848_), .A2(new_n672_), .A3(new_n555_), .A4(new_n886_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n903_), .A2(new_n904_), .A3(G190gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n903_), .B2(G190gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n902_), .B1(new_n905_), .B2(new_n906_), .ZN(G1351gat));
  INV_X1    g706(.A(new_n886_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n841_), .A2(new_n872_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n346_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT126), .B1(new_n910_), .B2(new_n342_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n342_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n909_), .A2(new_n913_), .A3(G197gat), .A4(new_n346_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n912_), .A3(new_n914_), .ZN(G1352gat));
  NOR4_X1   g714(.A1(new_n841_), .A2(new_n300_), .A3(new_n872_), .A4(new_n908_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n290_), .ZN(G1353gat));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919_));
  INV_X1    g718(.A(G211gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n873_), .A2(new_n626_), .A3(new_n886_), .A4(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n919_), .A2(new_n920_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n918_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n841_), .A2(new_n688_), .A3(new_n872_), .A4(new_n908_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n925_), .A2(new_n921_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n923_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n925_), .A2(KEYINPUT127), .A3(new_n921_), .A4(new_n927_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n924_), .A2(new_n926_), .A3(new_n928_), .ZN(G1354gat));
  AOI21_X1  g728(.A(G218gat), .B1(new_n909_), .B2(new_n671_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n672_), .A2(G218gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n909_), .B2(new_n931_), .ZN(G1355gat));
endmodule


