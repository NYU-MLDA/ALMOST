//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  OR2_X1    g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT25), .B(G183gat), .Z(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT26), .B(G190gat), .Z(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT78), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT79), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(new_n205_), .C1(new_n206_), .C2(new_n207_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n212_), .A3(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n209_), .A2(new_n214_), .A3(new_n216_), .A4(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n211_), .A2(new_n220_), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT81), .B(G176gat), .Z(new_n222_));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT22), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT22), .B1(new_n223_), .B2(new_n224_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n219_), .A2(KEYINPUT82), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT82), .B1(new_n219_), .B2(new_n228_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT21), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(KEYINPUT21), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n229_), .A2(new_n230_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT20), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n202_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G226gat), .A2(G233gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT88), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT19), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n219_), .A2(new_n228_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n219_), .A2(KEYINPUT82), .A3(new_n228_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n237_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n211_), .A2(new_n212_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT90), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n205_), .B(new_n251_), .C1(new_n253_), .C2(new_n207_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G169gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n222_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n221_), .A2(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259_));
  OR3_X1    g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n248_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n258_), .B2(new_n248_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n240_), .A2(new_n243_), .A3(new_n250_), .A4(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n248_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n239_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n237_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n266_), .B(new_n267_), .C1(new_n265_), .C2(new_n264_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n243_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n263_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT18), .B(G64gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G92gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n240_), .A2(new_n269_), .A3(new_n250_), .A4(new_n262_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n267_), .A2(KEYINPUT20), .A3(new_n264_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n243_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n275_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n282_), .A3(KEYINPUT27), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT1), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT84), .ZN(new_n286_));
  OR2_X1    g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n288_), .A3(KEYINPUT1), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(KEYINPUT85), .A3(new_n287_), .A4(new_n289_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n292_), .B(new_n293_), .C1(KEYINPUT1), .C2(new_n284_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT86), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n302_), .A2(KEYINPUT86), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n297_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(KEYINPUT3), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n295_), .A2(new_n302_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT87), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n307_), .A2(KEYINPUT87), .B1(new_n309_), .B2(new_n298_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .A4(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n301_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n314_));
  XOR2_X1   g113(.A(G78gat), .B(G106gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n248_), .B1(new_n313_), .B2(KEYINPUT29), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G22gat), .B(G50gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT28), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n317_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n325_), .A3(new_n316_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n263_), .A2(new_n281_), .A3(new_n270_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n281_), .B1(new_n263_), .B2(new_n270_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n283_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT98), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339_));
  INV_X1    g138(.A(G113gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G120gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n313_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT94), .B1(new_n345_), .B2(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n301_), .A2(new_n343_), .A3(new_n312_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n313_), .A2(new_n349_), .A3(new_n344_), .A4(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n346_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT93), .Z(new_n354_));
  AND2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n345_), .A2(new_n347_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(new_n354_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n355_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(new_n360_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n229_), .A2(new_n230_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT30), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n343_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(new_n343_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT31), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n373_), .A2(new_n343_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n374_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n371_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n370_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n331_), .A2(new_n283_), .A3(new_n336_), .A4(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n338_), .A2(new_n367_), .A3(new_n387_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n331_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n283_), .A2(new_n336_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n367_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n383_), .A2(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n271_), .B1(new_n396_), .B2(new_n281_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n280_), .A2(KEYINPUT32), .A3(new_n275_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n397_), .B(new_n398_), .C1(new_n364_), .C2(new_n366_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n361_), .B1(new_n362_), .B2(new_n354_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n354_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n346_), .A2(new_n348_), .A3(new_n401_), .A4(new_n351_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT96), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n403_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n400_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n263_), .A2(new_n270_), .A3(new_n281_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n276_), .A3(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT33), .B(new_n361_), .C1(new_n355_), .C2(new_n363_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n365_), .B2(new_n360_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n399_), .B(new_n331_), .C1(new_n408_), .C2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n394_), .A2(new_n395_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n390_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G148gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G176gat), .B(G204gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT70), .B(G120gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT68), .ZN(new_n424_));
  XOR2_X1   g223(.A(G85gat), .B(G92gat), .Z(new_n425_));
  INV_X1    g224(.A(KEYINPUT64), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT9), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT10), .B(G99gat), .Z(new_n431_));
  INV_X1    g230(.A(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n426_), .A2(new_n427_), .A3(G85gat), .A4(G92gat), .ZN(new_n434_));
  AND3_X1   g233(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT65), .B1(new_n435_), .B2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n448_));
  NAND3_X1  g247(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(new_n444_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n439_), .B1(new_n451_), .B2(new_n425_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n425_), .A2(new_n439_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n437_), .B2(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n438_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT67), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT67), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n438_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n460_));
  INV_X1    g259(.A(G57gat), .ZN(new_n461_));
  INV_X1    g260(.A(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G57gat), .A2(G64gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G71gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT66), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT66), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G71gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G78gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT66), .B(G71gat), .ZN(new_n473_));
  INV_X1    g272(.A(G78gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n463_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n466_), .A2(new_n472_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n473_), .A2(new_n474_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n468_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n465_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT12), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n459_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G230gat), .A2(G233gat), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT12), .B1(new_n455_), .B2(new_n482_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n481_), .B(new_n438_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n486_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n455_), .A2(new_n482_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n489_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n424_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n424_), .B1(new_n494_), .B2(new_n491_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n417_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n424_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n495_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  INV_X1    g306(.A(G50gat), .ZN(new_n508_));
  AND2_X1   g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n509_), .A2(new_n510_), .A3(G43gat), .ZN(new_n511_));
  INV_X1    g310(.A(G43gat), .ZN(new_n512_));
  INV_X1    g311(.A(G29gat), .ZN(new_n513_));
  INV_X1    g312(.A(G36gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n512_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n508_), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(G43gat), .B1(new_n509_), .B2(new_n510_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(G50gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G1gat), .B(G8gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(G1gat), .A2(G8gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT14), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G15gat), .A2(G22gat), .ZN(new_n526_));
  AND2_X1   g325(.A1(G15gat), .A2(G22gat), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n523_), .B(new_n525_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G8gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT74), .B1(new_n522_), .B2(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n519_), .A2(new_n520_), .A3(G50gat), .ZN(new_n534_));
  AOI21_X1  g333(.A(G50gat), .B1(new_n519_), .B2(new_n520_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n529_), .B(new_n523_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT74), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n518_), .A2(KEYINPUT15), .A3(new_n521_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT15), .B1(new_n518_), .B2(new_n521_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n532_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT76), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n540_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n522_), .A2(new_n532_), .A3(KEYINPUT75), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(new_n550_), .B2(new_n540_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n507_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n224_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(G197gat), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n548_), .A2(new_n549_), .B1(new_n533_), .B2(new_n539_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n540_), .A2(new_n543_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n545_), .ZN(new_n560_));
  OAI22_X1  g359(.A1(new_n558_), .A2(new_n544_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n507_), .A3(new_n555_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n506_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n415_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n541_), .A2(new_n542_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n459_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n438_), .B(new_n536_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n572_), .A2(new_n574_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G134gat), .ZN(new_n582_));
  INV_X1    g381(.A(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n576_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n459_), .B2(new_n568_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n585_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n578_), .B1(new_n588_), .B2(new_n575_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n567_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n593_));
  NOR4_X1   g392(.A1(new_n593_), .A2(new_n572_), .A3(new_n574_), .A4(new_n587_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT37), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n532_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n482_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT16), .B(G183gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G211gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n600_), .A2(KEYINPUT17), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT73), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(KEYINPUT17), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n590_), .A2(new_n595_), .A3(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n597_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n566_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(G1gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n393_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT99), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n612_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n596_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n566_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n367_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n619_), .A2(KEYINPUT99), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(KEYINPUT99), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT38), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n626_), .A3(new_n629_), .ZN(G1324gat));
  NAND4_X1  g429(.A1(new_n415_), .A2(new_n624_), .A3(new_n565_), .A4(new_n392_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G8gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G8gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n566_), .A2(new_n616_), .ZN(new_n635_));
  INV_X1    g434(.A(G8gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n392_), .A2(new_n636_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n633_), .A2(new_n634_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT100), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640_));
  OAI221_X1 g439(.A(new_n640_), .B1(new_n635_), .B2(new_n637_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n639_), .A2(KEYINPUT40), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT40), .B1(new_n639_), .B2(new_n641_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n625_), .B2(new_n395_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n635_), .A2(G15gat), .A3(new_n395_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n331_), .A2(G22gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT101), .Z(new_n650_));
  NAND2_X1  g449(.A1(new_n617_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G22gat), .B1(new_n625_), .B2(new_n331_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(KEYINPUT42), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(KEYINPUT42), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n651_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT102), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(new_n651_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(new_n596_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n565_), .A2(new_n623_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n660_), .B(new_n661_), .C1(new_n390_), .C2(new_n414_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n513_), .A3(new_n393_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n590_), .A2(new_n595_), .A3(new_n613_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n613_), .B1(new_n590_), .B2(new_n595_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n415_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n415_), .A2(new_n671_), .A3(KEYINPUT43), .A4(new_n667_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n661_), .B(KEYINPUT103), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT105), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .A4(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n393_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G29gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G29gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n663_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(new_n669_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n415_), .B2(new_n667_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(KEYINPUT43), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n666_), .B(new_n688_), .C1(new_n390_), .C2(new_n414_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n673_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n687_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n392_), .B(new_n680_), .C1(new_n691_), .C2(new_n675_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n662_), .A2(new_n514_), .A3(new_n392_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(KEYINPUT46), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  AND3_X1   g499(.A1(new_n662_), .A2(new_n512_), .A3(new_n387_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n387_), .B(new_n680_), .C1(new_n691_), .C2(new_n675_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G43gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n706_), .B(new_n701_), .C1(new_n702_), .C2(G43gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n662_), .B2(new_n391_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n677_), .A2(new_n391_), .A3(new_n680_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G50gat), .ZN(G1331gat));
  AOI211_X1 g510(.A(new_n563_), .B(new_n505_), .C1(new_n390_), .C2(new_n414_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n616_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n393_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT108), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n624_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n716_), .A2(new_n461_), .A3(new_n367_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1332gat));
  INV_X1    g517(.A(new_n716_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n462_), .B1(new_n719_), .B2(new_n392_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT48), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n713_), .A2(new_n462_), .A3(new_n392_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n716_), .B2(new_n395_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n713_), .A2(new_n467_), .A3(new_n387_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  NAND3_X1  g526(.A1(new_n713_), .A2(new_n474_), .A3(new_n391_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G78gat), .B1(new_n716_), .B2(new_n331_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(KEYINPUT50), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT50), .B1(new_n730_), .B2(new_n731_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n732_), .B2(new_n733_), .ZN(G1335gat));
  NOR3_X1   g533(.A1(new_n505_), .A2(new_n612_), .A3(new_n563_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n415_), .A2(new_n596_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(G85gat), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(new_n393_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n670_), .A2(new_n672_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n393_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(G85gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n736_), .B2(new_n392_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n392_), .A2(G92gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n739_), .B2(new_n745_), .ZN(G1337gat));
  INV_X1    g545(.A(G99gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n739_), .B2(new_n387_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n736_), .A2(new_n431_), .A3(new_n387_), .ZN(new_n749_));
  OAI22_X1  g548(.A1(new_n748_), .A2(new_n749_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n750_));
  NAND2_X1  g549(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT112), .Z(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(new_n754_));
  OAI221_X1 g553(.A(new_n752_), .B1(KEYINPUT111), .B2(KEYINPUT51), .C1(new_n748_), .C2(new_n749_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1338gat));
  NAND3_X1  g555(.A1(new_n736_), .A2(new_n432_), .A3(new_n391_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n670_), .A2(new_n391_), .A3(new_n672_), .A4(new_n735_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  NAND2_X1  g565(.A1(new_n501_), .A2(new_n495_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n558_), .A2(new_n545_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n559_), .A2(new_n560_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n556_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n561_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n556_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n767_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT55), .B1(new_n486_), .B2(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n491_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n485_), .A2(KEYINPUT55), .A3(new_n490_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n423_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n486_), .A2(KEYINPUT115), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n485_), .A2(new_n490_), .A3(KEYINPUT55), .A4(new_n780_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT116), .B(new_n775_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n483_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n783_));
  NOR4_X1   g582(.A1(new_n783_), .A2(new_n492_), .A3(new_n489_), .A4(new_n487_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n776_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n778_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n423_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n781_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n782_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n491_), .A2(new_n494_), .A3(new_n423_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n563_), .A2(KEYINPUT114), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT114), .B1(new_n563_), .B2(new_n792_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n774_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n596_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n799_));
  NOR2_X1   g598(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n788_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n779_), .A2(new_n781_), .A3(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n772_), .A2(new_n792_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n800_), .ZN(new_n808_));
  AND4_X1   g607(.A1(new_n787_), .A2(new_n786_), .A3(new_n781_), .A4(new_n801_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n801_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n799_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n806_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n807_), .A2(new_n814_), .A3(new_n667_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n788_), .A2(new_n789_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n775_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT56), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n795_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n596_), .B1(new_n819_), .B2(new_n773_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n815_), .B1(KEYINPUT57), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n798_), .B1(new_n821_), .B2(KEYINPUT120), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n797_), .B1(new_n796_), .B2(new_n596_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n815_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n612_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n496_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n416_), .B1(new_n501_), .B2(new_n495_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n564_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT113), .B1(new_n615_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n563_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n666_), .A2(new_n831_), .A3(new_n832_), .A4(new_n612_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n830_), .A2(KEYINPUT54), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT54), .B1(new_n830_), .B2(new_n833_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n826_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  AND4_X1   g637(.A1(new_n393_), .A2(new_n338_), .A3(new_n387_), .A4(new_n389_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(KEYINPUT119), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT119), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n837_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n820_), .A2(KEYINPUT57), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n823_), .A2(new_n844_), .A3(new_n815_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n623_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n836_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n839_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n843_), .A2(G113gat), .A3(new_n563_), .A4(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n340_), .B1(new_n849_), .B2(new_n564_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1340gat));
  OAI21_X1  g652(.A(new_n342_), .B1(new_n505_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT121), .B1(new_n342_), .B2(KEYINPUT60), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n849_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n854_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n843_), .A2(new_n506_), .A3(new_n850_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n860_), .B2(new_n342_), .ZN(G1341gat));
  NOR2_X1   g660(.A1(new_n849_), .A2(new_n623_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n843_), .A2(new_n612_), .A3(new_n850_), .ZN(new_n863_));
  MUX2_X1   g662(.A(new_n862_), .B(new_n863_), .S(G127gat), .Z(G1342gat));
  NOR2_X1   g663(.A1(new_n849_), .A2(new_n660_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n843_), .A2(new_n667_), .A3(new_n850_), .ZN(new_n866_));
  MUX2_X1   g665(.A(new_n865_), .B(new_n866_), .S(G134gat), .Z(G1343gat));
  AOI21_X1  g666(.A(new_n836_), .B1(new_n845_), .B2(new_n623_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n367_), .A3(new_n387_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n392_), .A2(new_n331_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n564_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n505_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g674(.A1(new_n871_), .A2(new_n623_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT61), .B(G155gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  NOR3_X1   g677(.A1(new_n871_), .A2(new_n583_), .A3(new_n666_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n869_), .A2(new_n596_), .A3(new_n870_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n583_), .B2(new_n880_), .ZN(G1347gat));
  AOI21_X1  g680(.A(new_n393_), .B1(new_n336_), .B2(new_n283_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n387_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n391_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n563_), .B(new_n884_), .C1(new_n826_), .C2(new_n836_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G169gat), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(KEYINPUT62), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n884_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n815_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n819_), .A2(new_n773_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n893_), .B2(new_n660_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n892_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n844_), .A3(new_n825_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n623_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n891_), .B1(new_n897_), .B2(new_n847_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n563_), .A2(new_n255_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT123), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n886_), .A2(new_n887_), .A3(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n890_), .A2(new_n901_), .A3(new_n903_), .ZN(G1348gat));
  OAI21_X1  g703(.A(new_n884_), .B1(new_n826_), .B2(new_n836_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n222_), .B1(new_n905_), .B2(new_n505_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n848_), .A2(KEYINPUT124), .A3(new_n331_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n868_), .B2(new_n391_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n883_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n907_), .A2(new_n909_), .A3(G176gat), .A4(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n906_), .B1(new_n505_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n906_), .B(KEYINPUT125), .C1(new_n505_), .C2(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1349gat));
  NAND4_X1  g715(.A1(new_n907_), .A2(new_n909_), .A3(new_n612_), .A4(new_n910_), .ZN(new_n917_));
  INV_X1    g716(.A(G183gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n253_), .B(new_n884_), .C1(new_n826_), .C2(new_n836_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n623_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n898_), .A2(KEYINPUT126), .A3(new_n612_), .A4(new_n253_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n919_), .A2(new_n922_), .A3(new_n923_), .A4(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n905_), .B2(new_n666_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n660_), .A2(new_n207_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n905_), .B2(new_n930_), .ZN(G1351gat));
  AND2_X1   g730(.A1(new_n848_), .A2(new_n882_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n387_), .A2(new_n331_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n563_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n506_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  AND2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  NOR4_X1   g740(.A1(new_n934_), .A2(new_n623_), .A3(new_n940_), .A4(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n935_), .A2(new_n612_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n940_), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n935_), .B2(new_n596_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n934_), .A2(new_n666_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(G218gat), .B2(new_n946_), .ZN(G1355gat));
endmodule


