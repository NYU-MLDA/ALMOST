//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G85gat), .B(G92gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n215_), .B(new_n217_), .C1(new_n216_), .C2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n212_), .A2(KEYINPUT64), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT7), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(KEYINPUT64), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n218_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n220_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n212_), .ZN(new_n228_));
  AOI211_X1 g027(.A(KEYINPUT8), .B(new_n218_), .C1(new_n228_), .C2(new_n223_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n209_), .B(new_n219_), .C1(new_n227_), .C2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G232gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT34), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT35), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n219_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n208_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n233_), .A2(new_n234_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT69), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(KEYINPUT67), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n230_), .A2(new_n246_), .A3(new_n235_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n245_), .A2(new_n247_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n242_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n244_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G134gat), .B(G162gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT68), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G190gat), .B(G218gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT36), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT70), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n256_), .A3(KEYINPUT71), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT37), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n254_), .A2(KEYINPUT36), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n244_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n263_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n266_), .A2(new_n267_), .B1(KEYINPUT37), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT65), .B(G71gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G78gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G57gat), .B(G64gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT11), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n272_), .A2(KEYINPUT11), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G15gat), .A2(G22gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G15gat), .A2(G22gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G1gat), .A2(G8gat), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n283_), .A2(new_n284_), .B1(KEYINPUT14), .B2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(new_n286_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n279_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT17), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G183gat), .B(G211gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G127gat), .B(G155gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n290_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(KEYINPUT17), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n270_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT75), .B1(new_n290_), .B2(new_n298_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n269_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n277_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n238_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n277_), .B(new_n219_), .C1(new_n227_), .C2(new_n229_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(KEYINPUT12), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT12), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n238_), .A2(new_n309_), .A3(new_n305_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G230gat), .A2(G233gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n307_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT66), .B(KEYINPUT5), .Z(new_n318_));
  XNOR2_X1  g117(.A(G120gat), .B(G148gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT13), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n304_), .A2(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT76), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(KEYINPUT76), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332_));
  XOR2_X1   g131(.A(G64gat), .B(G92gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT94), .Z(new_n339_));
  INV_X1    g138(.A(G176gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT84), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT23), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n345_), .B2(KEYINPUT23), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G183gat), .A3(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT85), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n353_), .A2(new_n350_), .A3(G183gat), .A4(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT95), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n360_));
  AOI211_X1 g159(.A(new_n360_), .B(new_n357_), .C1(new_n349_), .C2(new_n355_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n344_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT96), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT96), .B(new_n344_), .C1(new_n359_), .C2(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(G204gat), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  INV_X1    g169(.A(G204gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G197gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(G211gat), .A2(G218gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT21), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n370_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT92), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n373_), .A4(new_n377_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n374_), .A2(new_n375_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n371_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n376_), .B1(G197gat), .B2(G204gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n369_), .A2(new_n376_), .A3(new_n372_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n388_), .A2(KEYINPUT90), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT90), .B1(new_n388_), .B2(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n384_), .A2(new_n392_), .ZN(new_n393_));
  OR3_X1    g192(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n338_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n345_), .A2(KEYINPUT23), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n351_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G183gat), .ZN(new_n402_));
  INV_X1    g201(.A(G183gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT25), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(G190gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n398_), .A2(new_n400_), .A3(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT93), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n366_), .A2(new_n393_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT19), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n384_), .A2(new_n392_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT26), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G190gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n402_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(KEYINPUT81), .B2(new_n404_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n404_), .A2(KEYINPUT81), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT82), .B(G190gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(KEYINPUT26), .ZN(new_n423_));
  AND2_X1   g222(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n421_), .B(KEYINPUT26), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n419_), .B(new_n420_), .C1(new_n423_), .C2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n397_), .B1(new_n349_), .B2(new_n355_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n343_), .A2(new_n338_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n403_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n430_), .A2(KEYINPUT86), .B1(new_n400_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n343_), .A2(new_n433_), .A3(new_n338_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n428_), .A2(new_n429_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n412_), .B(new_n414_), .C1(new_n415_), .C2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n384_), .A2(new_n435_), .A3(new_n392_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n438_), .A2(KEYINPUT20), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n409_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(new_n393_), .ZN(new_n441_));
  AOI221_X4 g240(.A(new_n337_), .B1(new_n411_), .B2(new_n437_), .C1(new_n441_), .C2(new_n414_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n337_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n414_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n411_), .A2(new_n437_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n332_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G127gat), .B(G134gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G120gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G155gat), .A2(G162gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT87), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G155gat), .A3(G162gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461_));
  INV_X1    g260(.A(G141gat), .ZN(new_n462_));
  INV_X1    g261(.A(G148gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n460_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G141gat), .B(G148gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n454_), .A2(new_n456_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT1), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n454_), .A2(new_n456_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n452_), .B1(new_n477_), .B2(KEYINPUT1), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n473_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n451_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT88), .B1(new_n474_), .B2(new_n452_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(new_n459_), .A3(new_n470_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n476_), .A2(new_n478_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n482_), .B(new_n450_), .C1(new_n483_), .C2(new_n473_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n484_), .A3(KEYINPUT4), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n451_), .C1(new_n472_), .C2(new_n479_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT98), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT99), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n485_), .A2(KEYINPUT99), .A3(new_n487_), .A4(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n480_), .A2(new_n484_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n488_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G1gat), .B(G29gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(G85gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n493_), .A2(new_n502_), .A3(new_n494_), .A4(new_n497_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT103), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT103), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n507_), .A3(new_n503_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n414_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n439_), .B(new_n510_), .C1(new_n440_), .C2(new_n393_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n362_), .A2(new_n384_), .A3(new_n392_), .A4(new_n408_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n512_), .B(KEYINPUT20), .C1(new_n393_), .C2(new_n435_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n414_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n337_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n444_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT27), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n447_), .A2(new_n509_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n520_));
  OAI221_X1 g319(.A(new_n482_), .B1(new_n483_), .B2(new_n473_), .C1(new_n415_), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G228gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT28), .ZN(new_n523_));
  XOR2_X1   g322(.A(G22gat), .B(G50gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n521_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n415_), .A2(new_n520_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G78gat), .B(G106gat), .Z(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  OR2_X1    g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n529_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n519_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n444_), .A2(new_n445_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n337_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT100), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT33), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n505_), .A2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n491_), .A2(new_n492_), .B1(new_n496_), .B2(new_n488_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n541_), .A2(new_n502_), .A3(new_n494_), .A4(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n489_), .B1(new_n495_), .B2(KEYINPUT101), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(KEYINPUT101), .B2(new_n495_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n503_), .A3(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n536_), .A2(new_n543_), .A3(new_n517_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n515_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT102), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT102), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n515_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n444_), .A2(new_n549_), .A3(new_n445_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n548_), .B(new_n532_), .C1(new_n556_), .C2(new_n509_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G227gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n450_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G15gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT31), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n559_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563_));
  INV_X1    g362(.A(G43gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n435_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n562_), .B(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n534_), .A2(new_n557_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT104), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n534_), .A2(new_n557_), .A3(KEYINPUT104), .A4(new_n567_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n519_), .A2(new_n533_), .A3(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n208_), .B(KEYINPUT77), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n289_), .A2(new_n240_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n208_), .B(KEYINPUT77), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n289_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n577_), .B1(new_n581_), .B2(new_n576_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT78), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(KEYINPUT78), .B2(new_n582_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT79), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G169gat), .B(G197gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n586_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT80), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n586_), .B(new_n589_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT80), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n574_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n330_), .A2(new_n331_), .A3(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n509_), .A2(G1gat), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT107), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT106), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n259_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT105), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n574_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n574_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n509_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n328_), .A2(new_n302_), .A3(new_n591_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n600_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n602_), .A2(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n447_), .A2(new_n518_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n604_), .B(KEYINPUT105), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n572_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT106), .B(new_n620_), .C1(new_n621_), .C2(new_n571_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n619_), .B(new_n613_), .C1(new_n622_), .C2(new_n607_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT110), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT110), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n623_), .A2(new_n627_), .A3(new_n624_), .A4(G8gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT109), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n630_), .B(new_n624_), .C1(new_n623_), .C2(G8gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n623_), .A2(G8gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT109), .B1(new_n632_), .B2(KEYINPUT39), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n629_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n618_), .A2(G8gat), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n330_), .A2(new_n331_), .A3(new_n597_), .A4(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n617_), .B1(new_n634_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n636_), .B(KEYINPUT108), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n633_), .A2(new_n631_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT40), .B(new_n640_), .C1(new_n641_), .C2(new_n629_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(G1325gat));
  NAND2_X1  g442(.A1(new_n610_), .A2(new_n613_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G15gat), .B1(new_n644_), .B2(new_n567_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT41), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n598_), .A2(G15gat), .A3(new_n567_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(KEYINPUT41), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(G1326gat));
  OAI21_X1  g448(.A(G22gat), .B1(new_n644_), .B2(new_n532_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT42), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n532_), .A2(G22gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n598_), .B2(new_n652_), .ZN(G1327gat));
  NOR3_X1   g452(.A1(new_n606_), .A2(new_n302_), .A3(new_n327_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n597_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n611_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n574_), .A2(new_n658_), .A3(new_n269_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT111), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n574_), .A2(new_n269_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT43), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n574_), .A2(KEYINPUT111), .A3(new_n269_), .A4(new_n658_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n327_), .A2(new_n302_), .A3(new_n593_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT44), .B1(new_n665_), .B2(new_n666_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n509_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n657_), .B1(new_n669_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n655_), .A2(new_n671_), .A3(new_n619_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n655_), .A2(KEYINPUT45), .A3(new_n671_), .A4(new_n619_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n667_), .A2(new_n668_), .A3(new_n618_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n671_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(KEYINPUT112), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n680_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n665_), .A2(new_n666_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n666_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n619_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n676_), .B1(new_n687_), .B2(G36gat), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n681_), .A2(new_n690_), .ZN(G1329gat));
  INV_X1    g490(.A(new_n567_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n655_), .A2(new_n564_), .A3(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n692_), .A3(new_n686_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G43gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g495(.A(G50gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n655_), .A2(new_n697_), .A3(new_n533_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n667_), .A2(new_n668_), .A3(new_n532_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n697_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT114), .B(new_n698_), .C1(new_n699_), .C2(new_n697_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1331gat));
  AOI211_X1 g503(.A(new_n328_), .B(new_n591_), .C1(new_n621_), .C2(new_n571_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n304_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n611_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n592_), .A2(new_n595_), .A3(new_n302_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n328_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n610_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n611_), .A2(G57gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1332gat));
  OAI21_X1  g512(.A(G64gat), .B1(new_n710_), .B2(new_n618_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT48), .ZN(new_n715_));
  INV_X1    g514(.A(G64gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n716_), .A3(new_n619_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1333gat));
  INV_X1    g517(.A(G71gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n706_), .A2(new_n719_), .A3(new_n692_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G71gat), .B1(new_n710_), .B2(new_n567_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT49), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT49), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT115), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n720_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n710_), .B2(new_n532_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  INV_X1    g529(.A(G78gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n706_), .A2(new_n731_), .A3(new_n533_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1335gat));
  AND3_X1   g532(.A1(new_n705_), .A2(new_n303_), .A3(new_n620_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n611_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n328_), .A2(new_n302_), .A3(new_n591_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n665_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n665_), .B2(new_n737_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n611_), .A2(G85gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n735_), .B1(new_n740_), .B2(new_n741_), .ZN(G1336gat));
  AOI21_X1  g541(.A(G92gat), .B1(new_n734_), .B2(new_n619_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n619_), .A2(G92gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n740_), .B2(new_n744_), .ZN(G1337gat));
  NAND3_X1  g544(.A1(new_n734_), .A2(new_n214_), .A3(new_n692_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n738_), .A2(new_n739_), .A3(new_n567_), .ZN(new_n747_));
  INV_X1    g546(.A(G99gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n746_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n665_), .A2(new_n533_), .A3(new_n737_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(G106gat), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n734_), .A2(new_n213_), .A3(new_n533_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n755_), .A2(new_n756_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT53), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n755_), .A2(new_n756_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n758_), .A4(new_n757_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1339gat));
  NAND2_X1  g564(.A1(new_n268_), .A2(KEYINPUT37), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n264_), .A2(new_n265_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n264_), .A2(new_n265_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n308_), .A2(new_n315_), .A3(new_n310_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(KEYINPUT55), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n770_), .B2(KEYINPUT55), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n313_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(KEYINPUT55), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(new_n312_), .A3(new_n311_), .A4(new_n772_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n778_), .A3(new_n323_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n775_), .A2(new_n778_), .A3(KEYINPUT56), .A4(new_n323_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(KEYINPUT120), .A3(new_n780_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n325_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n581_), .A2(new_n577_), .A3(new_n576_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n577_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n589_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n784_), .A2(new_n785_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n769_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT121), .B1(new_n792_), .B2(new_n793_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n785_), .A2(new_n791_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(KEYINPUT58), .A4(new_n784_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n794_), .A2(new_n795_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n591_), .A2(new_n325_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n790_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n606_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n303_), .B1(new_n799_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n708_), .A2(KEYINPUT118), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n592_), .A2(new_n595_), .A3(new_n809_), .A4(new_n302_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n328_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n807_), .B1(new_n812_), .B2(new_n769_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n811_), .A2(new_n269_), .A3(KEYINPUT54), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n806_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n533_), .A2(new_n567_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n619_), .A2(new_n509_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n816_), .A2(new_n821_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n820_), .A2(G113gat), .A3(new_n596_), .A4(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n819_), .B2(new_n593_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1340gat));
  NAND3_X1  g625(.A1(new_n820_), .A2(new_n327_), .A3(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n816_), .A2(new_n817_), .ZN(new_n829_));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(KEYINPUT60), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n328_), .A2(KEYINPUT60), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n829_), .A2(KEYINPUT122), .A3(new_n818_), .A4(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835_));
  INV_X1    g634(.A(new_n833_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n819_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(new_n838_), .ZN(G1341gat));
  NAND4_X1  g638(.A1(new_n820_), .A2(G127gat), .A3(new_n302_), .A4(new_n822_), .ZN(new_n840_));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n819_), .B2(new_n303_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n769_), .A2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT123), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n820_), .A2(new_n822_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n819_), .B2(new_n606_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n532_), .A2(new_n692_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n806_), .B2(new_n815_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n818_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n593_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT124), .B(G141gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n854_), .B(new_n856_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n853_), .A2(new_n328_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n463_), .ZN(G1345gat));
  NOR2_X1   g658(.A1(new_n853_), .A2(new_n303_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n860_), .B(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(new_n853_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n864_), .A2(G162gat), .A3(new_n269_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G162gat), .B1(new_n864_), .B2(new_n620_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1347gat));
  XOR2_X1   g666(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n618_), .A2(new_n611_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n816_), .A2(new_n817_), .A3(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n593_), .ZN(new_n872_));
  INV_X1    g671(.A(G169gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n342_), .B2(new_n341_), .ZN(new_n875_));
  OAI211_X1 g674(.A(G169gat), .B(new_n868_), .C1(new_n871_), .C2(new_n593_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(G1348gat));
  NOR2_X1   g676(.A1(new_n871_), .A2(new_n328_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n340_), .ZN(G1349gat));
  NOR3_X1   g678(.A1(new_n871_), .A2(new_n303_), .A3(new_n405_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n829_), .A2(new_n302_), .A3(new_n870_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n403_), .B2(new_n881_), .ZN(G1350gat));
  OAI21_X1  g681(.A(G190gat), .B1(new_n871_), .B2(new_n769_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n620_), .A2(new_n406_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n871_), .B2(new_n884_), .ZN(G1351gat));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n816_), .A2(new_n886_), .A3(new_n850_), .A4(new_n870_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n803_), .B(KEYINPUT57), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n794_), .A2(new_n795_), .A3(new_n798_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n302_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n813_), .A2(new_n814_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n850_), .B(new_n870_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT126), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n887_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G197gat), .B1(new_n894_), .B2(new_n591_), .ZN(new_n895_));
  INV_X1    g694(.A(G197gat), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n896_), .B(new_n593_), .C1(new_n887_), .C2(new_n893_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n327_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G204gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n371_), .A3(new_n327_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1353gat));
  OR2_X1    g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n894_), .B2(new_n302_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT63), .B(G211gat), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n303_), .B(new_n905_), .C1(new_n887_), .C2(new_n893_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1354gat));
  NAND2_X1  g706(.A1(new_n894_), .A2(new_n620_), .ZN(new_n908_));
  INV_X1    g707(.A(G218gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n769_), .A2(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT127), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n908_), .A2(new_n909_), .B1(new_n894_), .B2(new_n911_), .ZN(G1355gat));
endmodule


