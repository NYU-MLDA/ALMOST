//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202_));
  AND2_X1   g001(.A1(G127gat), .A2(G134gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G127gat), .ZN(new_n206_));
  INV_X1    g005(.A(G134gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G127gat), .A2(G134gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT82), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G113gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n205_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n213_));
  INV_X1    g012(.A(G120gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n203_), .A2(new_n204_), .A3(new_n202_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT82), .B1(new_n208_), .B2(new_n209_), .ZN(new_n217_));
  OAI21_X1  g016(.A(G113gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n205_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n219_));
  AOI21_X1  g018(.A(G120gat), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G155gat), .ZN(new_n221_));
  INV_X1    g020(.A(G162gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT83), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT83), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(G155gat), .B2(G162gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT84), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n223_), .A2(new_n225_), .A3(KEYINPUT84), .A4(new_n226_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT3), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT2), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n229_), .A2(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(KEYINPUT1), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(G155gat), .A3(G162gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n236_), .A2(new_n223_), .A3(new_n225_), .A4(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n231_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n233_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n215_), .A2(new_n220_), .B1(new_n235_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n214_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n229_), .A2(new_n230_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n232_), .A2(new_n234_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n218_), .A2(G120gat), .A3(new_n219_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n244_), .A2(new_n247_), .A3(new_n248_), .A4(new_n241_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n248_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n251_), .B(new_n252_), .C1(new_n235_), .C2(new_n242_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT93), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n243_), .A2(new_n249_), .A3(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G85gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n257_), .A3(new_n263_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(G176gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n268_), .A2(new_n269_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT23), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT80), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n278_), .A3(KEYINPUT23), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT81), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n275_), .B2(KEYINPUT23), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n282_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n277_), .A2(new_n279_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n274_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT25), .B(G183gat), .Z(new_n287_));
  INV_X1    g086(.A(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT26), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT77), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G190gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n294_), .A2(KEYINPUT76), .A3(KEYINPUT77), .A4(G190gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n287_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n275_), .B(KEYINPUT23), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n298_));
  INV_X1    g097(.A(G169gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n269_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT24), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n272_), .A2(new_n273_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n297_), .B(new_n303_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n286_), .B1(new_n296_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n251_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(new_n251_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G43gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT31), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n314_), .B(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G71gat), .B(G99gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT30), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G227gat), .A2(G233gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n318_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G78gat), .B(G106gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT88), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT89), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT29), .B1(new_n235_), .B2(new_n242_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT21), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(G204gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(G204gat), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n332_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G211gat), .B(G218gat), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n331_), .A2(G197gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT21), .B1(new_n336_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n332_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT21), .A3(new_n338_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(G233gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n329_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n329_), .B2(new_n345_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n328_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n352_), .A3(new_n327_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n235_), .A2(new_n242_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G22gat), .B(G50gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n361_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n366_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n364_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n328_), .B(KEYINPUT90), .C1(new_n353_), .C2(new_n354_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n359_), .A2(new_n368_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n326_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n368_), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT91), .B(new_n326_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n357_), .A4(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT98), .ZN(new_n381_));
  XOR2_X1   g180(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n382_));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n301_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n270_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n277_), .A2(new_n279_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n281_), .A2(new_n283_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n287_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n292_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n297_), .B1(G183gat), .B2(G190gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n274_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n345_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n388_), .A2(new_n307_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n297_), .A2(new_n303_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n295_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n294_), .A2(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n289_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT76), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n403_), .B1(new_n406_), .B2(new_n291_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n401_), .B(new_n402_), .C1(new_n407_), .C2(new_n287_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n342_), .A2(new_n344_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n286_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT19), .ZN(new_n412_));
  AND4_X1   g211(.A1(KEYINPUT20), .A2(new_n400_), .A3(new_n410_), .A4(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n310_), .B2(new_n345_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n398_), .A3(new_n396_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n387_), .B1(new_n413_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n310_), .A2(new_n345_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(KEYINPUT20), .A3(new_n416_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n412_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n400_), .A2(new_n410_), .A3(KEYINPUT20), .A4(new_n412_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n386_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n399_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n396_), .A2(KEYINPUT96), .A3(new_n398_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n409_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n421_), .B1(new_n431_), .B2(new_n415_), .ZN(new_n432_));
  AND4_X1   g231(.A1(KEYINPUT20), .A2(new_n400_), .A3(new_n410_), .A4(new_n421_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n386_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT27), .A3(new_n418_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n380_), .A2(new_n381_), .A3(new_n427_), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n427_), .A2(new_n435_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n373_), .A2(new_n379_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT98), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n267_), .B(new_n324_), .C1(new_n436_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n266_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n266_), .B2(new_n442_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n256_), .A2(KEYINPUT33), .A3(new_n257_), .A4(new_n263_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n250_), .A2(new_n254_), .A3(new_n253_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n243_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n264_), .A3(new_n448_), .ZN(new_n449_));
  AND4_X1   g248(.A1(new_n418_), .A2(new_n446_), .A3(new_n424_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n422_), .A2(new_n423_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n265_), .A2(new_n266_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT32), .B(new_n387_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n445_), .A2(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT97), .B1(new_n455_), .B2(new_n438_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n437_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n267_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n438_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n266_), .A2(new_n442_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT95), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n418_), .A2(new_n449_), .A3(new_n424_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n266_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n446_), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n453_), .A2(new_n454_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n380_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n456_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n440_), .B1(new_n469_), .B2(new_n324_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G230gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G85gat), .B(G92gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT6), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT64), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT64), .B1(new_n477_), .B2(new_n479_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n474_), .B(new_n475_), .C1(new_n482_), .C2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n477_), .A2(new_n479_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n474_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT8), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(G85gat), .A3(G92gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n473_), .B2(new_n491_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n482_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n490_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G71gat), .B(G78gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(KEYINPUT11), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n500_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT67), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n499_), .A2(new_n512_), .A3(KEYINPUT12), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT12), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n486_), .A2(new_n489_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n507_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n507_), .ZN(new_n517_));
  AND4_X1   g316(.A1(new_n472_), .A2(new_n513_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G176gat), .B(G204gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G120gat), .B(G148gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n499_), .A2(new_n510_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT66), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n526_), .A2(new_n517_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n519_), .B(new_n524_), .C1(new_n527_), .C2(new_n472_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n524_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n472_), .B1(new_n526_), .B2(new_n517_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(new_n518_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(KEYINPUT69), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT69), .B1(new_n528_), .B2(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n471_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT13), .A3(new_n532_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT73), .B(G1gat), .Z(new_n539_));
  INV_X1    g338(.A(G8gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT14), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G1gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G8gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n543_), .B(G1gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n540_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(G43gat), .ZN(new_n550_));
  INV_X1    g349(.A(G29gat), .ZN(new_n551_));
  INV_X1    g350(.A(G36gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(G50gat), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(G50gat), .B1(new_n556_), .B2(new_n557_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n549_), .A2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n546_), .B(new_n548_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(KEYINPUT75), .A3(new_n563_), .ZN(new_n564_));
  OR3_X1    g363(.A1(new_n549_), .A2(KEYINPUT75), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  INV_X1    g368(.A(G50gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n557_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n555_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n569_), .B1(new_n572_), .B2(new_n558_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n558_), .A3(new_n569_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(KEYINPUT15), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT15), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n573_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n546_), .A2(new_n548_), .A3(new_n576_), .A4(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n562_), .A2(new_n566_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n568_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n299_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n334_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n585_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n470_), .A2(new_n538_), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G134gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n222_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n576_), .A2(new_n579_), .A3(new_n499_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n515_), .A2(new_n561_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n598_), .A2(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n595_), .A2(new_n605_), .A3(new_n600_), .A4(new_n601_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n594_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n592_), .A2(new_n593_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT71), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT72), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n604_), .A2(KEYINPUT72), .A3(new_n606_), .A4(new_n609_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n607_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI211_X1 g415(.A(KEYINPUT37), .B(new_n607_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n549_), .B(new_n619_), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n507_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n512_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n620_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n620_), .A2(new_n629_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(KEYINPUT17), .A3(new_n631_), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n618_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n589_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n267_), .A3(new_n539_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT99), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n638_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n634_), .A2(new_n614_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n589_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n458_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n641_), .A3(new_n645_), .ZN(G1324gat));
  NAND3_X1  g445(.A1(new_n636_), .A2(new_n540_), .A3(new_n437_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n437_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G8gat), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT39), .B(new_n540_), .C1(new_n643_), .C2(new_n437_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT100), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n654_), .B(new_n647_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n643_), .B2(new_n323_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n636_), .A2(new_n658_), .A3(new_n323_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n643_), .B2(new_n438_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT101), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n636_), .A2(new_n663_), .A3(new_n438_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n634_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n614_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n589_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n551_), .A3(new_n267_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n618_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n470_), .A2(KEYINPUT43), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n469_), .A2(new_n324_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n440_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(KEYINPUT103), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n670_), .A2(KEYINPUT37), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n614_), .A2(new_n615_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(KEYINPUT104), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n470_), .A2(KEYINPUT103), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n470_), .B2(KEYINPUT103), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n467_), .B1(new_n466_), .B2(new_n380_), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT97), .B(new_n438_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n323_), .B1(new_n698_), .B2(new_n459_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n699_), .B2(new_n440_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n694_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n678_), .B1(new_n693_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n535_), .A2(new_n537_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n588_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n634_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n707_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n708_), .A2(new_n709_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n676_), .B1(new_n703_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n678_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT105), .B1(new_n701_), .B2(KEYINPUT43), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n692_), .B(new_n715_), .C1(new_n694_), .C2(new_n700_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n676_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n710_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n458_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n673_), .B1(new_n720_), .B2(new_n551_), .ZN(G1328gat));
  XNOR2_X1  g520(.A(new_n437_), .B(KEYINPUT107), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n672_), .A2(new_n552_), .A3(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT45), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n457_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n552_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT46), .B(new_n724_), .C1(new_n725_), .C2(new_n552_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  AOI211_X1 g529(.A(new_n550_), .B(new_n324_), .C1(new_n712_), .C2(new_n719_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n672_), .A2(new_n323_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n550_), .A2(KEYINPUT108), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n550_), .A2(KEYINPUT108), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT47), .B1(new_n731_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n712_), .A2(new_n719_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(G43gat), .A3(new_n323_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n735_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1330gat));
  NAND3_X1  g541(.A1(new_n672_), .A2(new_n570_), .A3(new_n438_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n380_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n570_), .ZN(G1331gat));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n470_), .A2(new_n705_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT109), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT109), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n538_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n635_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n751_), .B2(new_n458_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT110), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n538_), .A3(new_n642_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n754_), .A2(new_n746_), .A3(new_n458_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1332gat));
  INV_X1    g555(.A(new_n722_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G64gat), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT48), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n757_), .A2(G64gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n751_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n754_), .B2(new_n324_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n324_), .A2(G71gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n751_), .B2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n754_), .B2(new_n380_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n380_), .A2(G78gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n751_), .B2(new_n768_), .ZN(G1335gat));
  AND4_X1   g568(.A1(new_n538_), .A2(new_n748_), .A3(new_n671_), .A4(new_n749_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n267_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT111), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n705_), .A2(new_n669_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n538_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n703_), .A2(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n267_), .A2(G85gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1336gat));
  NAND3_X1  g576(.A1(new_n775_), .A2(G92gat), .A3(new_n722_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n770_), .A2(new_n437_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(G92gat), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT112), .ZN(G1337gat));
  NAND3_X1  g580(.A1(new_n770_), .A2(new_n495_), .A3(new_n323_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n774_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n717_), .A2(new_n323_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G99gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G99gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT51), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n782_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1338gat));
  NAND3_X1  g591(.A1(new_n717_), .A2(new_n438_), .A3(new_n783_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(G106gat), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n770_), .A2(new_n496_), .A3(new_n438_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT114), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n770_), .A2(new_n800_), .A3(new_n496_), .A4(new_n438_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n797_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n796_), .A2(new_n805_), .A3(new_n797_), .A4(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  NAND2_X1  g606(.A1(new_n436_), .A2(new_n439_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n323_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n528_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n472_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n516_), .A2(new_n517_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n513_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n518_), .B1(new_n816_), .B2(KEYINPUT55), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NOR4_X1   g617(.A1(new_n814_), .A2(new_n815_), .A3(new_n818_), .A4(new_n813_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n529_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT115), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n816_), .A2(KEYINPUT55), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n519_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n819_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n524_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n822_), .A2(new_n823_), .B1(new_n827_), .B2(KEYINPUT56), .ZN(new_n828_));
  AOI211_X1 g627(.A(KEYINPUT116), .B(new_n821_), .C1(new_n820_), .C2(KEYINPUT115), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n812_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n585_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n562_), .A2(new_n567_), .A3(new_n580_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n835_), .A3(new_n585_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n536_), .A2(new_n586_), .A3(new_n532_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n830_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n839_), .B2(new_n670_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n841_), .B(new_n614_), .C1(new_n830_), .C2(new_n838_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n827_), .B2(KEYINPUT56), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n820_), .A2(new_n845_), .A3(new_n821_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n846_), .C1(new_n821_), .C2(new_n820_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n837_), .A2(new_n586_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n528_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n847_), .A2(new_n848_), .A3(KEYINPUT58), .A4(new_n528_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n618_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n669_), .B1(new_n843_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n635_), .A2(new_n588_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT54), .B1(new_n855_), .B2(new_n538_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n704_), .A2(new_n635_), .A3(new_n857_), .A4(new_n588_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n267_), .B(new_n810_), .C1(new_n854_), .C2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n705_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(KEYINPUT59), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n851_), .A2(new_n618_), .A3(new_n852_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n859_), .B1(new_n866_), .B2(new_n669_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n267_), .A4(new_n810_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n864_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n588_), .A2(new_n211_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n863_), .B1(new_n870_), .B2(new_n871_), .ZN(G1340gat));
  NAND3_X1  g671(.A1(new_n864_), .A2(new_n869_), .A3(new_n538_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n214_), .B1(new_n704_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n862_), .B(new_n875_), .C1(KEYINPUT60), .C2(new_n214_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(KEYINPUT119), .A3(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n634_), .B2(KEYINPUT120), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n870_), .B(new_n882_), .C1(KEYINPUT120), .C2(G127gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n206_), .B1(new_n861_), .B2(new_n634_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n862_), .B2(new_n614_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n677_), .A2(new_n207_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n870_), .B2(new_n887_), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n843_), .A2(new_n853_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n860_), .B1(new_n889_), .B2(new_n634_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(new_n323_), .A3(new_n380_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n267_), .A3(new_n757_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n588_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT121), .B(G141gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  AND2_X1   g694(.A1(new_n891_), .A2(new_n267_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n538_), .A3(new_n757_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n669_), .A3(new_n757_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT122), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n899_), .B(new_n901_), .ZN(G1346gat));
  NOR3_X1   g701(.A1(new_n892_), .A2(new_n222_), .A3(new_n687_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n896_), .A2(new_n614_), .A3(new_n757_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n222_), .B2(new_n904_), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n890_), .A2(new_n438_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n757_), .A2(new_n267_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n323_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT123), .Z(new_n909_));
  NAND3_X1  g708(.A1(new_n906_), .A2(new_n705_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT124), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n906_), .A2(new_n912_), .A3(new_n705_), .A4(new_n909_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(G169gat), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n906_), .A2(new_n909_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(new_n705_), .A3(new_n268_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n911_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n913_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(G1348gat));
  NOR2_X1   g719(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n538_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n922_), .B2(new_n921_), .ZN(G1349gat));
  NAND2_X1  g724(.A1(new_n917_), .A2(new_n669_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G183gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n287_), .B2(new_n926_), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n917_), .A2(new_n292_), .A3(new_n614_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n917_), .A2(new_n618_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n288_), .ZN(G1351gat));
  NAND2_X1  g730(.A1(new_n891_), .A2(new_n907_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n588_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n334_), .ZN(G1352gat));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  OAI22_X1  g734(.A1(new_n932_), .A2(new_n704_), .B1(new_n935_), .B2(G204gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(G204gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT127), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n936_), .B(new_n938_), .ZN(G1353gat));
  INV_X1    g738(.A(new_n932_), .ZN(new_n940_));
  AOI211_X1 g739(.A(KEYINPUT63), .B(G211gat), .C1(new_n940_), .C2(new_n669_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT63), .B(G211gat), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n932_), .A2(new_n634_), .A3(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1354gat));
  AND3_X1   g743(.A1(new_n940_), .A2(G218gat), .A3(new_n618_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G218gat), .B1(new_n940_), .B2(new_n614_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1355gat));
endmodule


