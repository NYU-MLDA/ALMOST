//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n208_), .B(new_n211_), .Z(new_n212_));
  NAND2_X1  g011(.A1(G229gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(new_n208_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n208_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n211_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n215_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G113gat), .B(G141gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G169gat), .B(G197gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT84), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G113gat), .B(G120gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT31), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT82), .B(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(G169gat), .B2(G176gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT23), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n233_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT80), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT24), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(G183gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G190gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n251_), .C1(new_n252_), .C2(new_n248_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n237_), .B(KEYINPUT81), .ZN(new_n257_));
  INV_X1    g056(.A(new_n239_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n241_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265_));
  INV_X1    g064(.A(G43gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n264_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(G15gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT30), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n268_), .B(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n230_), .B1(new_n273_), .B2(KEYINPUT85), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(KEYINPUT85), .B2(new_n273_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n273_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n230_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G197gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT91), .B1(new_n280_), .B2(G204gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(G204gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n280_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT21), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n280_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT92), .B1(new_n280_), .B2(G204gat), .ZN(new_n288_));
  OAI22_X1  g087(.A1(new_n287_), .A2(new_n288_), .B1(new_n280_), .B2(G204gat), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n285_), .B(new_n286_), .C1(new_n289_), .C2(KEYINPUT21), .ZN(new_n290_));
  INV_X1    g089(.A(new_n286_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(KEYINPUT21), .A3(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT88), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT88), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n304_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n303_), .B(new_n305_), .C1(new_n306_), .C2(KEYINPUT2), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT89), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n301_), .A2(new_n307_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n298_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n297_), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT86), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(KEYINPUT1), .B2(new_n297_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n314_), .A2(new_n315_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n306_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n313_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n294_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n326_), .A2(G228gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(G228gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G78gat), .ZN(new_n330_));
  INV_X1    g129(.A(G106gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n324_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n323_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT28), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n322_), .A2(new_n336_), .A3(new_n323_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G22gat), .B(G50gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n333_), .B1(new_n343_), .B2(KEYINPUT93), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT93), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(KEYINPUT93), .A3(new_n333_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n293_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n233_), .B1(new_n259_), .B2(new_n234_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n240_), .B1(new_n254_), .B2(new_n242_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n252_), .A2(new_n251_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n247_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n293_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n365_), .A2(KEYINPUT20), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n262_), .A2(new_n263_), .A3(new_n293_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n361_), .A2(new_n364_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n294_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n358_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n355_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT100), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT100), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n375_), .B(new_n355_), .C1(new_n367_), .C2(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n365_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(KEYINPUT20), .A3(new_n358_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n365_), .A2(new_n377_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n359_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n358_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n374_), .A2(new_n376_), .B1(new_n354_), .B2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G1gat), .B(G29gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  INV_X1    g188(.A(new_n321_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n229_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n310_), .B(KEYINPUT89), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n390_), .B(new_n391_), .C1(new_n392_), .C2(new_n298_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n229_), .B1(new_n313_), .B2(new_n321_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT95), .B(new_n229_), .C1(new_n313_), .C2(new_n321_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT97), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  INV_X1    g200(.A(new_n399_), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n401_), .B(new_n402_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n396_), .A2(KEYINPUT4), .A3(new_n397_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n394_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n399_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n389_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n402_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n389_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n411_), .B(new_n412_), .C1(new_n400_), .C2(new_n403_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n409_), .B1(new_n413_), .B2(KEYINPUT101), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT101), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n398_), .A2(new_n399_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n401_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n398_), .A2(KEYINPUT97), .A3(new_n399_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n419_), .B2(new_n412_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n384_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT98), .B1(new_n413_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n399_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n424_));
  AOI211_X1 g223(.A(new_n412_), .B(new_n424_), .C1(new_n410_), .C2(new_n399_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n383_), .A2(new_n353_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n353_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n381_), .A2(new_n427_), .A3(new_n382_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT98), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n419_), .A2(new_n430_), .A3(KEYINPUT33), .A4(new_n412_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n413_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n423_), .A2(new_n429_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n349_), .B1(new_n421_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n428_), .A2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n427_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n347_), .A2(new_n437_), .A3(new_n440_), .A4(new_n348_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n441_), .A2(new_n414_), .A3(new_n420_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n279_), .B1(new_n435_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n414_), .A2(new_n420_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n279_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n440_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n349_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n225_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT10), .B(G99gat), .Z(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT64), .B(G106gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT6), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT67), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(KEYINPUT67), .B2(new_n461_), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT66), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(G92gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT65), .B(G85gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT9), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n464_), .A2(new_n471_), .A3(KEYINPUT68), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT68), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n474_));
  OR2_X1    g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n461_), .A2(KEYINPUT67), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT9), .ZN(new_n480_));
  AND2_X1   g279(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT66), .B(G92gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n473_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n460_), .B1(new_n472_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G85gat), .B(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n455_), .A2(new_n457_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n331_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n488_), .B(new_n490_), .C1(new_n491_), .C2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT70), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT70), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(new_n490_), .C1(new_n491_), .C2(new_n496_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(KEYINPUT8), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(KEYINPUT70), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G78gat), .Z(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n487_), .A2(new_n501_), .A3(new_n503_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT71), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n495_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n489_), .B1(new_n516_), .B2(new_n458_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n499_), .B1(new_n517_), .B2(new_n488_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n503_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n521_), .A2(KEYINPUT71), .A3(new_n487_), .A4(new_n510_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n487_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n510_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n513_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT68), .B1(new_n464_), .B2(new_n471_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n479_), .A2(new_n485_), .A3(new_n473_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n459_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n532_), .B2(new_n510_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n534_), .B(new_n524_), .C1(new_n520_), .C2(new_n531_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n533_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n528_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G176gat), .B(G204gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT73), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n528_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n546_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT75), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n539_), .A2(new_n545_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n557_), .A3(KEYINPUT13), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n510_), .B(new_n208_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n571_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n573_), .B2(new_n565_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n532_), .A2(new_n211_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n523_), .A2(new_n216_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT76), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT34), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT35), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n579_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n577_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n582_), .A2(new_n583_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n577_), .A2(new_n578_), .A3(new_n588_), .A4(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT36), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n596_), .A3(new_n589_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n594_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT77), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT37), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n602_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n576_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n450_), .A2(new_n562_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n203_), .A3(new_n445_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n598_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n225_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n576_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n562_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT103), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n445_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n616_), .A2(KEYINPUT104), .A3(G1gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT104), .B1(new_n616_), .B2(G1gat), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n609_), .B1(new_n617_), .B2(new_n618_), .ZN(G1324gat));
  NAND3_X1  g418(.A1(new_n606_), .A2(new_n204_), .A3(new_n447_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT105), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n610_), .A2(new_n614_), .A3(new_n621_), .A4(new_n447_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(G8gat), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n610_), .A2(new_n614_), .A3(new_n447_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT105), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n624_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT40), .B(new_n620_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1325gat));
  INV_X1    g432(.A(new_n279_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n606_), .A2(new_n270_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n615_), .A2(new_n634_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n636_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(new_n636_), .B2(G15gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(G1326gat));
  INV_X1    g438(.A(G22gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n349_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT106), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n606_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n615_), .A2(new_n349_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G22gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT42), .B(new_n640_), .C1(new_n615_), .C2(new_n349_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(G1327gat));
  INV_X1    g447(.A(new_n562_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(new_n225_), .A3(new_n612_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n443_), .A2(new_n449_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n603_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n604_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n658_), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n660_), .B(new_n652_), .C1(new_n443_), .C2(new_n449_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n650_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT44), .B(new_n650_), .C1(new_n659_), .C2(new_n661_), .ZN(new_n665_));
  AND4_X1   g464(.A1(G29gat), .A2(new_n664_), .A3(new_n445_), .A4(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n598_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n612_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n562_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n450_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n445_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n666_), .A2(new_n672_), .ZN(G1328gat));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n447_), .A3(new_n665_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G36gat), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n671_), .A2(new_n676_), .A3(new_n447_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT45), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n675_), .A2(new_n678_), .A3(KEYINPUT46), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1329gat));
  NAND4_X1  g482(.A1(new_n664_), .A2(G43gat), .A3(new_n634_), .A4(new_n665_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n266_), .B1(new_n670_), .B2(new_n279_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1330gat));
  AND4_X1   g487(.A1(G50gat), .A2(new_n664_), .A3(new_n349_), .A4(new_n665_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G50gat), .B1(new_n671_), .B2(new_n349_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n562_), .A2(new_n611_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(new_n605_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n445_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n610_), .A2(new_n612_), .A3(new_n692_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n445_), .B2(KEYINPUT109), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(KEYINPUT109), .B2(new_n698_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n697_), .B2(new_n700_), .ZN(G1332gat));
  INV_X1    g500(.A(G64gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n697_), .B2(new_n447_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n695_), .A2(new_n702_), .A3(new_n447_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n697_), .B2(new_n634_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT49), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n279_), .A2(G71gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT111), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n695_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n697_), .B2(new_n349_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT50), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n349_), .A2(new_n715_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT112), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n695_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1335gat));
  AND2_X1   g520(.A1(new_n694_), .A2(new_n668_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n445_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n659_), .A2(new_n661_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n693_), .A2(new_n612_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n444_), .A2(new_n483_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(G1336gat));
  AOI21_X1  g527(.A(G92gat), .B1(new_n722_), .B2(new_n447_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n484_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n726_), .B2(new_n730_), .ZN(G1337gat));
  AND3_X1   g530(.A1(new_n722_), .A2(new_n634_), .A3(new_n451_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n634_), .A3(new_n725_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G99gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n734_), .B(new_n735_), .Z(G1338gat));
  XNOR2_X1  g535(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n349_), .B(new_n725_), .C1(new_n659_), .C2(new_n661_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G106gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n738_), .A3(G106gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n722_), .A2(new_n349_), .A3(new_n452_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n737_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n742_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n744_), .B(new_n737_), .C1(new_n746_), .C2(new_n740_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1339gat));
  INV_X1    g548(.A(KEYINPUT122), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n611_), .A2(G113gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n634_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT55), .B(new_n533_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n535_), .A2(new_n537_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n513_), .A2(new_n522_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n527_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT12), .B1(new_n532_), .B2(new_n510_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n536_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n533_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n538_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n756_), .A2(new_n759_), .A3(new_n762_), .A4(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n545_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n212_), .A2(new_n213_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n224_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n213_), .B1(new_n220_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n217_), .A2(KEYINPUT119), .A3(new_n219_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n221_), .A2(new_n773_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n778_), .A2(new_n779_), .A3(KEYINPUT120), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT120), .B1(new_n778_), .B2(new_n779_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n547_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n771_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n771_), .A2(new_n783_), .A3(KEYINPUT58), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n658_), .A3(new_n787_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n766_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n766_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT117), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n767_), .A2(KEYINPUT117), .A3(new_n768_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n611_), .A2(new_n547_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT118), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n769_), .A2(new_n797_), .A3(new_n770_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n793_), .B1(new_n790_), .B2(KEYINPUT117), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n552_), .A2(new_n557_), .A3(new_n782_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n796_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n667_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n788_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n798_), .A2(new_n800_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n802_), .B1(new_n808_), .B2(KEYINPUT118), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n598_), .B1(new_n809_), .B2(new_n801_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT57), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n612_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n561_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT13), .B1(new_n552_), .B2(new_n557_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n605_), .B(new_n225_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT115), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n562_), .A2(new_n817_), .A3(new_n225_), .A4(new_n605_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n818_), .A3(KEYINPUT54), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n753_), .B1(new_n812_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n753_), .C1(new_n812_), .C2(new_n823_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n786_), .A2(new_n658_), .A3(new_n787_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n810_), .B2(KEYINPUT57), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n805_), .A2(new_n806_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n576_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n816_), .A2(new_n818_), .A3(KEYINPUT54), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT54), .B1(new_n816_), .B2(new_n818_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT121), .A3(new_n825_), .A4(new_n753_), .ZN(new_n837_));
  AOI221_X4 g636(.A(new_n751_), .B1(KEYINPUT59), .B2(new_n824_), .C1(new_n828_), .C2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n752_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n611_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n750_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n840_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n828_), .A2(new_n837_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT122), .B(new_n842_), .C1(new_n845_), .C2(new_n751_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n562_), .B1(new_n824_), .B2(KEYINPUT59), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n843_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n562_), .A2(KEYINPUT60), .ZN(new_n851_));
  MUX2_X1   g650(.A(KEYINPUT60), .B(new_n851_), .S(new_n848_), .Z(new_n852_));
  NAND2_X1  g651(.A1(new_n839_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT123), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n649_), .B1(new_n839_), .B2(new_n825_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n828_), .B2(new_n837_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n856_), .B(new_n853_), .C1(new_n858_), .C2(new_n848_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(G1341gat));
  AOI21_X1  g659(.A(G127gat), .B1(new_n839_), .B2(new_n612_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n845_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n576_), .A2(KEYINPUT124), .ZN(new_n863_));
  MUX2_X1   g662(.A(KEYINPUT124), .B(new_n863_), .S(G127gat), .Z(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n862_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n824_), .B2(new_n667_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT125), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n660_), .A2(new_n866_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n862_), .B2(new_n869_), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n812_), .A2(new_n823_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n871_), .A2(new_n444_), .A3(new_n441_), .A4(new_n634_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n611_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT126), .B(G141gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n649_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n612_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n881_), .A3(new_n598_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n872_), .A2(new_n658_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1347gat));
  INV_X1    g683(.A(new_n349_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n446_), .A2(new_n885_), .A3(new_n447_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n871_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n611_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G169gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT127), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n891_), .A3(G169gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(KEYINPUT62), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n888_), .B2(G169gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  INV_X1    g694(.A(new_n888_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n232_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n897_), .ZN(G1348gat));
  NAND2_X1  g697(.A1(new_n887_), .A2(new_n649_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n245_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n231_), .B2(new_n899_), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n887_), .A2(new_n612_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n252_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n235_), .B2(new_n902_), .ZN(G1350gat));
  INV_X1    g703(.A(new_n887_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G190gat), .B1(new_n905_), .B2(new_n660_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n887_), .A2(new_n251_), .A3(new_n598_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1351gat));
  NAND3_X1  g707(.A1(new_n279_), .A2(new_n349_), .A3(new_n447_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n871_), .A2(new_n445_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n611_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n649_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n612_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  AND2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n915_), .B2(new_n916_), .ZN(G1354gat));
  INV_X1    g718(.A(G218gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n910_), .A2(new_n920_), .A3(new_n598_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n910_), .A2(new_n658_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n920_), .ZN(G1355gat));
endmodule


