//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT3), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n206_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n213_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n207_), .A3(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n220_), .B(KEYINPUT28), .Z(new_n221_));
  XOR2_X1   g020(.A(G197gat), .B(G204gat), .Z(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT21), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT21), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G211gat), .B(G218gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(KEYINPUT29), .B2(new_n219_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n221_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G78gat), .B(G106gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT98), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G228gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G22gat), .B(G50gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n231_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(G183gat), .ZN(new_n239_));
  INV_X1    g038(.A(G190gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT23), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT89), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT90), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT88), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT24), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT91), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n252_), .A3(new_n249_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n239_), .A3(KEYINPUT25), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT25), .B(G183gat), .Z(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n254_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT87), .B1(new_n258_), .B2(G190gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT26), .B(G190gat), .Z(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT87), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n257_), .A2(new_n261_), .B1(new_n248_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n251_), .A2(new_n253_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT92), .B1(new_n267_), .B2(KEYINPUT22), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT22), .B(G169gat), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n266_), .B(new_n268_), .C1(new_n269_), .C2(KEYINPUT92), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n241_), .A2(new_n244_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n239_), .A2(new_n240_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n273_), .A3(new_n262_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276_));
  INV_X1    g075(.A(G43gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n275_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT95), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G113gat), .B(G120gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n281_), .A2(KEYINPUT95), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(KEYINPUT95), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n283_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT96), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n288_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n280_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n280_), .A2(new_n294_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT94), .B(G15gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT93), .B(KEYINPUT30), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT97), .B(KEYINPUT31), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n295_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n238_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n295_), .A2(new_n296_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n303_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n231_), .B(new_n237_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n295_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT104), .ZN(new_n314_));
  INV_X1    g113(.A(new_n219_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(KEYINPUT4), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n316_), .A2(KEYINPUT102), .B1(new_n289_), .B2(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n294_), .A2(new_n219_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT102), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n322_), .B2(KEYINPUT4), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT103), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n314_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n329_));
  OAI211_X1 g128(.A(KEYINPUT104), .B(new_n325_), .C1(new_n329_), .C2(new_n317_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT106), .B1(new_n322_), .B2(new_n325_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT106), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n318_), .A2(new_n321_), .A3(new_n332_), .A4(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G1gat), .B(G29gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT105), .B(KEYINPUT0), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n327_), .A2(new_n340_), .A3(new_n330_), .A4(new_n334_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n313_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n249_), .A2(new_n271_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n256_), .A2(new_n260_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n248_), .A2(new_n263_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT99), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT99), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n269_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n262_), .B1(new_n353_), .B2(G176gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n246_), .B2(new_n272_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n228_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(KEYINPUT20), .B(new_n356_), .C1(new_n275_), .C2(new_n228_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT100), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n355_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n349_), .A2(new_n351_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n229_), .B(new_n366_), .C1(new_n367_), .C2(new_n345_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT20), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n229_), .B1(new_n265_), .B2(new_n274_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n359_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT100), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n357_), .A2(new_n374_), .A3(new_n359_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n361_), .A2(new_n365_), .A3(new_n373_), .A4(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT101), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n361_), .A2(new_n375_), .A3(new_n373_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n365_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n360_), .A2(KEYINPUT100), .B1(new_n371_), .B2(new_n372_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(KEYINPUT101), .A3(new_n365_), .A4(new_n375_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n378_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT109), .B(KEYINPUT27), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n371_), .A2(new_n372_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n357_), .A2(new_n359_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n376_), .B(KEYINPUT27), .C1(new_n365_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n344_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n343_), .A2(KEYINPUT107), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT33), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n343_), .A2(KEYINPUT107), .A3(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n318_), .A2(new_n321_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n340_), .B1(new_n397_), .B2(new_n325_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n378_), .A2(new_n399_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n394_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT108), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n382_), .A2(new_n403_), .A3(new_n375_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT108), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(new_n404_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n304_), .A2(new_n305_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n238_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n392_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n418_));
  NAND2_X1  g217(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G99gat), .A2(G106gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT6), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT10), .B(G99gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT64), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT65), .B(G85gat), .Z(new_n426_));
  INV_X1    g225(.A(KEYINPUT9), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n428_), .A2(G92gat), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT66), .ZN(new_n431_));
  OAI221_X1 g230(.A(new_n422_), .B1(new_n425_), .B2(G106gat), .C1(new_n429_), .C2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n433_));
  INV_X1    g232(.A(G99gat), .ZN(new_n434_));
  INV_X1    g233(.A(G106gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  XOR2_X1   g238(.A(G85gat), .B(G92gat), .Z(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n437_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT68), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n445_), .A3(new_n437_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n421_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .A4(new_n447_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n444_), .A2(new_n446_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n439_), .B1(new_n453_), .B2(new_n440_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n441_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AOI211_X1 g255(.A(KEYINPUT69), .B(new_n439_), .C1(new_n453_), .C2(new_n440_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n432_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G71gat), .B(G78gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G64gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(KEYINPUT11), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT70), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n461_), .A2(KEYINPUT70), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(KEYINPUT70), .ZN(new_n466_));
  INV_X1    g265(.A(new_n463_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n420_), .B1(new_n458_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G230gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n458_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n446_), .A2(new_n452_), .A3(new_n450_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n445_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n440_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT8), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT69), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n454_), .A2(new_n455_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n441_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n464_), .A2(new_n468_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n432_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n458_), .A2(new_n469_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT71), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n472_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n481_), .A2(KEYINPUT71), .A3(new_n482_), .A4(new_n432_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G120gat), .B(G148gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n484_), .A2(new_n490_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n418_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n484_), .A2(new_n490_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(KEYINPUT13), .A3(new_n497_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G169gat), .B(G197gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  NAND2_X1  g308(.A1(G1gat), .A2(G8gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT14), .ZN(new_n511_));
  INV_X1    g310(.A(G15gat), .ZN(new_n512_));
  INV_X1    g311(.A(G22gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(G15gat), .A2(G22gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n511_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT80), .Z(new_n517_));
  XOR2_X1   g316(.A(G1gat), .B(G8gat), .Z(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(new_n518_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT15), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529_));
  INV_X1    g328(.A(new_n526_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n525_), .A2(new_n530_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n522_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n521_), .A2(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n521_), .A2(new_n527_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(new_n536_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n509_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n536_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n537_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n509_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n504_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n417_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n534_), .A2(new_n458_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n481_), .A2(new_n432_), .A3(new_n527_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT78), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n553_), .A2(new_n563_), .A3(new_n554_), .A4(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT76), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT77), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n562_), .A2(new_n564_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(KEYINPUT37), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n570_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT79), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n565_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n562_), .A2(KEYINPUT79), .A3(new_n564_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n577_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n576_), .B1(new_n582_), .B2(KEYINPUT37), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT81), .ZN(new_n584_));
  INV_X1    g383(.A(G231gat), .ZN(new_n585_));
  INV_X1    g384(.A(G233gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n482_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n464_), .A2(new_n589_), .A3(new_n468_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n588_), .A2(new_n590_), .A3(new_n521_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n521_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n584_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n590_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n589_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n522_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n590_), .A3(new_n521_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT81), .A3(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT16), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n602_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n597_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT83), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n596_), .A2(new_n597_), .A3(KEYINPUT83), .A4(new_n606_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n583_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n552_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n342_), .A2(new_n343_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n613_), .A2(G1gat), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n417_), .A2(new_n582_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n551_), .A2(new_n611_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n615_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n617_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n622_), .A3(new_n623_), .ZN(G1324gat));
  AND2_X1   g423(.A1(new_n386_), .A2(new_n390_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n613_), .A2(G8gat), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(new_n391_), .A3(new_n620_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n628_), .A3(G8gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(G8gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n621_), .B2(new_n414_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n414_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n512_), .ZN(new_n639_));
  OAI22_X1  g438(.A1(new_n636_), .A2(new_n637_), .B1(new_n613_), .B2(new_n639_), .ZN(G1326gat));
  XNOR2_X1  g439(.A(new_n238_), .B(KEYINPUT110), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n621_), .B2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(KEYINPUT42), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(KEYINPUT42), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(G22gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT111), .Z(new_n646_));
  OAI22_X1  g445(.A1(new_n643_), .A2(new_n644_), .B1(new_n613_), .B2(new_n646_), .ZN(G1327gat));
  NAND2_X1  g446(.A1(new_n565_), .A2(new_n579_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n581_), .A3(new_n570_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n575_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n611_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n552_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n614_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n551_), .A2(new_n651_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n415_), .B1(new_n402_), .B2(new_n412_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n657_), .B(new_n583_), .C1(new_n658_), .C2(new_n392_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n625_), .A2(new_n615_), .A3(new_n313_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n400_), .B1(new_n393_), .B2(KEYINPUT33), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n411_), .B1(new_n662_), .B2(new_n396_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n663_), .B2(new_n415_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n657_), .B1(new_n664_), .B2(new_n583_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT44), .B(new_n656_), .C1(new_n660_), .C2(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(G29gat), .A3(new_n614_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n660_), .A2(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n656_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n655_), .B1(new_n667_), .B2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT37), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n577_), .A2(new_n675_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n650_), .A2(new_n675_), .B1(new_n571_), .B2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n417_), .B2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n670_), .B1(new_n678_), .B2(new_n659_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n625_), .B1(new_n679_), .B2(KEYINPUT44), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n674_), .B1(new_n680_), .B2(new_n671_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n625_), .A2(G36gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT45), .B1(new_n653_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n552_), .A2(new_n685_), .A3(new_n652_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n673_), .B1(new_n681_), .B2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n679_), .A2(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n666_), .A2(new_n391_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G36gat), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(KEYINPUT46), .A3(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n689_), .A2(new_n693_), .ZN(G1329gat));
  OAI21_X1  g493(.A(new_n277_), .B1(new_n653_), .B2(new_n414_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n666_), .A2(G43gat), .A3(new_n638_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n690_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT47), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n695_), .C1(new_n696_), .C2(new_n690_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1330gat));
  INV_X1    g500(.A(G50gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n653_), .B2(new_n641_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n666_), .A2(G50gat), .A3(new_n310_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n690_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n707_), .B(new_n703_), .C1(new_n704_), .C2(new_n690_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1331gat));
  NAND4_X1  g508(.A1(new_n619_), .A2(new_n651_), .A3(new_n549_), .A4(new_n504_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n615_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n504_), .A2(new_n549_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n417_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n612_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n615_), .A2(G57gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n710_), .B2(new_n625_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(KEYINPUT48), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(KEYINPUT48), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n625_), .A2(G64gat), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT113), .Z(new_n721_));
  OAI22_X1  g520(.A1(new_n718_), .A2(new_n719_), .B1(new_n714_), .B2(new_n721_), .ZN(G1333gat));
  OR3_X1    g521(.A1(new_n714_), .A2(G71gat), .A3(new_n414_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G71gat), .B1(new_n710_), .B2(new_n414_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n725_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(G1334gat));
  OR3_X1    g527(.A1(new_n714_), .A2(G78gat), .A3(new_n641_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G78gat), .B1(new_n710_), .B2(new_n641_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT50), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT50), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n713_), .A2(new_n652_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n614_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n712_), .A2(new_n651_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n669_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n615_), .A2(new_n426_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n736_), .B1(new_n741_), .B2(new_n742_), .ZN(G1336gat));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n735_), .A2(new_n744_), .A3(new_n391_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n669_), .A2(new_n625_), .A3(new_n740_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n744_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT116), .ZN(G1337gat));
  NOR3_X1   g547(.A1(new_n734_), .A2(new_n425_), .A3(new_n414_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n638_), .B(new_n739_), .C1(new_n660_), .C2(new_n665_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(G99gat), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n751_), .B(new_n753_), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n735_), .A2(new_n435_), .A3(new_n310_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n310_), .B(new_n739_), .C1(new_n660_), .C2(new_n665_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n755_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  AOI21_X1  g563(.A(new_n482_), .B1(new_n481_), .B2(new_n432_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n474_), .B(new_n483_), .C1(new_n765_), .C2(new_n420_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n488_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT120), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n484_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n483_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n470_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n772_), .A2(KEYINPUT55), .A3(new_n472_), .A4(new_n474_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n766_), .A2(new_n774_), .A3(new_n488_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n768_), .A2(new_n770_), .A3(new_n773_), .A4(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n495_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n495_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(KEYINPUT121), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n495_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(KEYINPUT121), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n542_), .A2(new_n537_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n535_), .A2(new_n536_), .A3(new_n543_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n509_), .A3(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n547_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n497_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n782_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT122), .B1(new_n779_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n780_), .A2(new_n781_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n495_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n787_), .B1(new_n778_), .B2(KEYINPUT121), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n792_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(new_n583_), .A3(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n549_), .A2(new_n498_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n786_), .B1(new_n499_), .B2(new_n498_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n650_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n807_), .B(new_n582_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n651_), .B1(new_n801_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n611_), .A2(new_n548_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n583_), .A2(new_n812_), .A3(KEYINPUT118), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT118), .B1(new_n583_), .B2(new_n812_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n814_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n811_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n677_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT119), .B1(new_n823_), .B2(KEYINPUT54), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n813_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n810_), .A2(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n615_), .A2(new_n391_), .A3(new_n306_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n548_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n805_), .A2(new_n650_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n807_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n650_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n583_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n792_), .B(KEYINPUT58), .C1(new_n796_), .C2(new_n797_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n835_), .B(new_n836_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n611_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n818_), .A2(new_n819_), .A3(new_n814_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n813_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n829_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT59), .B(new_n829_), .C1(new_n810_), .C2(new_n827_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n833_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT123), .A3(new_n846_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n548_), .A2(G113gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT124), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n832_), .B1(new_n852_), .B2(new_n854_), .ZN(G1340gat));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  INV_X1    g655(.A(new_n504_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n831_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n856_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n850_), .B2(new_n846_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g660(.A(G127gat), .B1(new_n831_), .B2(new_n651_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n651_), .A2(G127gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n852_), .B2(new_n863_), .ZN(G1342gat));
  AOI21_X1  g663(.A(G134gat), .B1(new_n831_), .B2(new_n582_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n583_), .A2(G134gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n852_), .B2(new_n866_), .ZN(G1343gat));
  INV_X1    g666(.A(new_n312_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n844_), .A2(new_n614_), .A3(new_n625_), .A4(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n549_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n202_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n857_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n203_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n611_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n874_), .B(new_n876_), .ZN(G1346gat));
  INV_X1    g676(.A(G162gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n869_), .A2(new_n878_), .A3(new_n677_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n869_), .B2(new_n650_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT125), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(new_n878_), .C1(new_n869_), .C2(new_n650_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n881_), .B2(new_n883_), .ZN(G1347gat));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n625_), .A2(new_n614_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n638_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n641_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n549_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n885_), .B1(new_n828_), .B2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n844_), .A2(KEYINPUT126), .A3(new_n890_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(G169gat), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n892_), .A2(new_n893_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n844_), .A2(new_n269_), .A3(new_n890_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(G1348gat));
  NOR2_X1   g698(.A1(new_n828_), .A2(new_n889_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G176gat), .B1(new_n900_), .B2(new_n504_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n828_), .A2(new_n310_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n887_), .A2(new_n266_), .A3(new_n857_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n651_), .A3(new_n888_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n651_), .A2(new_n256_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n905_), .A2(new_n239_), .B1(new_n900_), .B2(new_n906_), .ZN(G1350gat));
  NOR2_X1   g706(.A1(new_n650_), .A2(new_n260_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n900_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n583_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n240_), .ZN(G1351gat));
  AOI21_X1  g711(.A(new_n312_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n548_), .A3(new_n886_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n504_), .A3(new_n886_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918_));
  INV_X1    g717(.A(G211gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n913_), .A2(new_n886_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n918_), .B(new_n919_), .C1(new_n920_), .C2(new_n611_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n919_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n611_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n913_), .A2(new_n886_), .A3(new_n922_), .A4(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n920_), .B2(new_n677_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n650_), .A2(G218gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n920_), .B2(new_n930_), .ZN(G1355gat));
endmodule


