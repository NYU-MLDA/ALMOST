//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT23), .A3(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT22), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT84), .A3(G169gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n216_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT82), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n222_), .A2(KEYINPUT24), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(KEYINPUT82), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n206_), .A2(new_n210_), .A3(new_n207_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .A4(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT25), .B(G183gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT81), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n221_), .B1(new_n230_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT30), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT30), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n240_), .B(new_n221_), .C1(new_n230_), .C2(new_n237_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n203_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n203_), .A3(new_n241_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G15gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n202_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n248_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n244_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(new_n242_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n249_), .A3(KEYINPUT87), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G127gat), .B(G134gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT85), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(KEYINPUT85), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n252_), .A2(new_n256_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n202_), .B(new_n268_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT19), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT94), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n229_), .A2(new_n209_), .B1(G169gat), .B2(G176gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n217_), .A2(G169gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n214_), .A2(KEYINPUT22), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT95), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT95), .B1(new_n276_), .B2(new_n277_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n216_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n233_), .A2(new_n225_), .A3(new_n223_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n208_), .A2(new_n211_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n275_), .A2(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G197gat), .B(G204gat), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT21), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT21), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G211gat), .ZN(new_n289_));
  INV_X1    g088(.A(G218gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT91), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT91), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n295_), .A3(new_n292_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n285_), .A2(new_n288_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n299_));
  OAI211_X1 g098(.A(KEYINPUT21), .B(new_n284_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n300_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n238_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n274_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n238_), .A2(new_n303_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n275_), .A2(new_n280_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n281_), .A2(new_n282_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n272_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n306_), .A2(new_n309_), .A3(KEYINPUT20), .A4(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G36gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT97), .B(G8gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n315_), .B(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n305_), .A2(new_n311_), .A3(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n306_), .A2(KEYINPUT20), .A3(new_n309_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n320_), .A2(KEYINPUT100), .A3(new_n272_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT100), .B1(new_n320_), .B2(new_n272_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n302_), .A2(new_n304_), .A3(new_n274_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(KEYINPUT27), .B(new_n319_), .C1(new_n324_), .C2(new_n318_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT90), .B(G228gat), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G233gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(KEYINPUT92), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329_));
  INV_X1    g128(.A(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G148gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n335_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n334_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n340_), .A2(new_n339_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n333_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n353_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n345_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n329_), .B1(new_n344_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n328_), .B1(new_n357_), .B2(new_n301_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n327_), .A2(KEYINPUT92), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n345_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n352_), .A2(new_n353_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n352_), .A2(new_n353_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT29), .B1(new_n364_), .B2(new_n343_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n365_), .B2(new_n303_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n358_), .B1(new_n366_), .B2(new_n328_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT93), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT28), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n344_), .A2(new_n356_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(KEYINPUT29), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n344_), .A2(new_n356_), .A3(new_n329_), .A4(new_n372_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n370_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n367_), .A2(new_n369_), .A3(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n358_), .B(new_n368_), .C1(new_n366_), .C2(new_n328_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n359_), .B1(new_n357_), .B2(new_n301_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n328_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n375_), .A2(new_n376_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n368_), .A4(new_n358_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n367_), .A2(new_n369_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n378_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n318_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n311_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n307_), .A2(new_n308_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n303_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n301_), .B(new_n221_), .C1(new_n230_), .C2(new_n237_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n273_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n319_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT102), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT102), .ZN(new_n401_));
  AOI211_X1 g200(.A(new_n401_), .B(KEYINPUT27), .C1(new_n397_), .C2(new_n319_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n325_), .B(new_n389_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT103), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n305_), .A2(new_n311_), .A3(new_n318_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n318_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n401_), .B1(new_n408_), .B2(KEYINPUT27), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n398_), .A2(KEYINPUT102), .A3(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n411_), .A2(KEYINPUT103), .A3(new_n325_), .A4(new_n389_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n270_), .B1(new_n405_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G85gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(G1gat), .B(G29gat), .Z(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n262_), .A2(new_n263_), .B1(new_n344_), .B2(new_n356_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(KEYINPUT4), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n374_), .A2(new_n261_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT4), .B1(new_n422_), .B2(new_n419_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n422_), .A2(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n418_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n417_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n418_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n374_), .A2(new_n261_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n264_), .A2(new_n374_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n429_), .B1(new_n433_), .B2(new_n420_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n417_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n426_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n428_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n267_), .A2(new_n269_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n411_), .A2(new_n438_), .A3(new_n325_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n389_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n318_), .A2(KEYINPUT32), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n443_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n322_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n320_), .A2(KEYINPUT100), .A3(new_n272_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n443_), .B1(new_n447_), .B2(new_n323_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n437_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT101), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n435_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n421_), .A2(new_n423_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(KEYINPUT99), .A3(new_n418_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT99), .B1(new_n452_), .B2(new_n418_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT98), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n436_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n436_), .A2(new_n458_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n456_), .B(new_n408_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT101), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n437_), .A2(new_n448_), .A3(new_n462_), .A4(new_n444_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n450_), .A2(new_n461_), .A3(new_n389_), .A4(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n413_), .A2(new_n438_), .B1(new_n442_), .B2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT71), .B(G43gat), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G50gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(G29gat), .B(G36gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT71), .B(G43gat), .ZN(new_n469_));
  INV_X1    g268(.A(G50gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n467_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n468_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n474_), .B(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n474_), .A2(new_n481_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n467_), .A2(new_n471_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n468_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n467_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT15), .A3(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n483_), .B1(new_n491_), .B2(new_n481_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  MUX2_X1   g292(.A(new_n482_), .B(new_n492_), .S(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(KEYINPUT80), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G113gat), .B(G141gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G169gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G197gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT10), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT10), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G99gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(G106gat), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT6), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT65), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n507_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(KEYINPUT65), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(KEYINPUT6), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n506_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n505_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517_));
  OR2_X1    g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n520_), .A2(KEYINPUT64), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n524_));
  AND2_X1   g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT9), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n527_), .B2(new_n521_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n516_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT66), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n516_), .B(new_n531_), .C1(new_n523_), .C2(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n513_), .A2(new_n514_), .A3(new_n506_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n506_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n534_), .B(new_n535_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n525_), .A2(new_n526_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n538_), .A2(KEYINPUT8), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT8), .B1(new_n538_), .B2(new_n539_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G78gat), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n533_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT12), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n551_), .A2(KEYINPUT12), .ZN(new_n555_));
  INV_X1    g354(.A(new_n541_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n538_), .A2(KEYINPUT8), .A3(new_n539_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n532_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT64), .B1(new_n520_), .B2(new_n522_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n527_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n531_), .B1(new_n561_), .B2(new_n516_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n556_), .B(new_n557_), .C1(new_n558_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n549_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n555_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n555_), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n549_), .B(new_n566_), .C1(new_n533_), .C2(new_n542_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n553_), .B(new_n554_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n564_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT67), .A3(new_n550_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n563_), .A2(KEYINPUT67), .A3(new_n564_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n554_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT70), .B(G120gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n568_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT13), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(KEYINPUT13), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n465_), .A2(new_n500_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT34), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT35), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n485_), .A2(new_n490_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n533_), .B2(new_n542_), .ZN(new_n594_));
  OAI211_X1 g393(.A(KEYINPUT35), .B(new_n591_), .C1(new_n594_), .C2(KEYINPUT72), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n563_), .A2(new_n474_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n594_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n563_), .A2(new_n491_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT72), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n474_), .B2(new_n563_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n591_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n592_), .B1(new_n598_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT75), .B(G190gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n605_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n605_), .B2(new_n614_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n589_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n598_), .A2(new_n604_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n612_), .B(new_n611_), .C1(new_n618_), .C2(new_n592_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n605_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT37), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n549_), .B(new_n481_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT79), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n628_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n627_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n622_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n588_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n588_), .A2(KEYINPUT104), .A3(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n476_), .A3(new_n437_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n615_), .A2(new_n616_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n640_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n588_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n438_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n653_), .ZN(G1324gat));
  NAND2_X1  g453(.A1(new_n411_), .A2(new_n325_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G8gat), .B1(new_n652_), .B2(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT105), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(KEYINPUT105), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(KEYINPUT39), .A3(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n647_), .A2(new_n477_), .A3(new_n655_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(KEYINPUT105), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(new_n666_), .A3(new_n661_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(KEYINPUT40), .A3(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  NOR3_X1   g471(.A1(new_n646_), .A2(G15gat), .A3(new_n270_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT107), .Z(new_n674_));
  OAI21_X1  g473(.A(G15gat), .B1(new_n652_), .B2(new_n270_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT41), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1326gat));
  OR3_X1    g476(.A1(new_n646_), .A2(G22gat), .A3(new_n389_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G22gat), .B1(new_n652_), .B2(new_n389_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT108), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n640_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n587_), .A2(new_n685_), .A3(new_n500_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n622_), .B2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n615_), .A2(new_n616_), .A3(new_n589_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT37), .B1(new_n619_), .B2(new_n620_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n465_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n692_), .B2(KEYINPUT109), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n405_), .A2(new_n412_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n442_), .A2(new_n464_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n694_), .B1(new_n698_), .B2(new_n622_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n686_), .B1(new_n693_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n686_), .C1(new_n693_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n438_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n650_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n465_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n686_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n708_), .A2(G29gat), .A3(new_n438_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n702_), .A2(new_n655_), .A3(new_n703_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n702_), .A2(KEYINPUT110), .A3(new_n655_), .A4(new_n703_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(G36gat), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n713_), .A2(KEYINPUT111), .A3(G36gat), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n708_), .A2(G36gat), .A3(new_n656_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT45), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(KEYINPUT46), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  OAI21_X1  g525(.A(G43gat), .B1(new_n704_), .B2(new_n270_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n439_), .A2(new_n203_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n708_), .B2(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n704_), .B2(new_n389_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n441_), .A2(new_n470_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n708_), .B2(new_n732_), .ZN(G1331gat));
  INV_X1    g532(.A(new_n586_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n584_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n500_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n698_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n641_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n437_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G57gat), .B1(new_n438_), .B2(KEYINPUT112), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n651_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(KEYINPUT112), .A2(G57gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n741_), .B1(new_n742_), .B2(new_n745_), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n743_), .B2(new_n656_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT48), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n656_), .A2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n739_), .B2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n743_), .B2(new_n270_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n270_), .A2(G71gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n739_), .B2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n743_), .B2(new_n389_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n389_), .A2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n739_), .B2(new_n757_), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n737_), .A2(new_n640_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n465_), .A3(new_n706_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n437_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n759_), .B(KEYINPUT113), .Z(new_n762_));
  NOR2_X1   g561(.A1(new_n693_), .A2(new_n699_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n762_), .A2(new_n438_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n655_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n762_), .A2(new_n656_), .A3(new_n763_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G92gat), .ZN(G1337gat));
  AOI21_X1  g567(.A(new_n270_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n760_), .A2(new_n769_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n762_), .A2(new_n270_), .A3(new_n763_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n501_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g572(.A(G106gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n760_), .A2(new_n774_), .A3(new_n441_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n762_), .A2(new_n763_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n441_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(G106gat), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT52), .B(new_n774_), .C1(new_n777_), .C2(new_n441_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n775_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  MUX2_X1   g581(.A(new_n492_), .B(new_n482_), .S(new_n493_), .Z(new_n783_));
  MUX2_X1   g582(.A(new_n494_), .B(new_n783_), .S(new_n499_), .Z(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT118), .B1(new_n568_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n550_), .A2(new_n552_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n569_), .A2(new_n566_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n563_), .A2(new_n564_), .A3(new_n555_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT55), .A4(new_n554_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n786_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n553_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n553_), .B(KEYINPUT117), .C1(new_n565_), .C2(new_n567_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n572_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT116), .B1(new_n568_), .B2(new_n785_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n568_), .A2(KEYINPUT116), .A3(new_n785_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n793_), .B(new_n798_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n579_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n568_), .A2(new_n785_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n568_), .A2(KEYINPUT116), .A3(new_n785_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(KEYINPUT119), .A3(new_n793_), .A4(new_n798_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n798_), .B1(new_n800_), .B2(new_n799_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n786_), .A2(new_n792_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n802_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n579_), .ZN(new_n814_));
  AND4_X1   g613(.A1(KEYINPUT56), .A2(new_n813_), .A3(new_n814_), .A4(new_n809_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n580_), .B(new_n784_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n813_), .A2(new_n814_), .A3(new_n809_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n809_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n580_), .A4(new_n784_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(new_n622_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n736_), .A2(new_n580_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n583_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n828_), .A2(new_n784_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n706_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT57), .B(new_n706_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n825_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n640_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT114), .B1(new_n736_), .B2(new_n640_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n692_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n685_), .A2(new_n839_), .A3(new_n500_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n735_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT115), .B1(new_n838_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n838_), .A2(new_n841_), .A3(KEYINPUT115), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n836_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n838_), .A2(new_n841_), .A3(KEYINPUT115), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(KEYINPUT54), .A3(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n835_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n413_), .A2(new_n437_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT120), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n736_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n835_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n834_), .A2(KEYINPUT121), .A3(new_n640_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n849_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n852_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n853_), .A2(KEYINPUT59), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n500_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n855_), .B1(new_n864_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g664(.A(G120gat), .B1(new_n863_), .B2(new_n735_), .ZN(new_n866_));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n735_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n854_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n867_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g669(.A(G127gat), .B1(new_n854_), .B2(new_n685_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n861_), .A2(G127gat), .A3(new_n862_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n685_), .ZN(G1342gat));
  AOI21_X1  g672(.A(G134gat), .B1(new_n854_), .B2(new_n650_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n863_), .A2(new_n692_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n656_), .A2(new_n437_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n850_), .A2(new_n270_), .A3(new_n441_), .A4(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n848_), .B1(new_n834_), .B2(new_n640_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n882_), .A2(new_n439_), .A3(new_n389_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT122), .B1(new_n883_), .B2(new_n878_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n736_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G141gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n879_), .A2(new_n880_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n882_), .A2(new_n439_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(KEYINPUT122), .A3(new_n441_), .A4(new_n878_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n330_), .A3(new_n736_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n886_), .A2(new_n891_), .ZN(G1344gat));
  OAI21_X1  g691(.A(new_n587_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G148gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n331_), .A3(new_n587_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1345gat));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n890_), .B2(new_n685_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n897_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n640_), .B(new_n899_), .C1(new_n887_), .C2(new_n889_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n890_), .B2(new_n650_), .ZN(new_n902_));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  AOI211_X1 g702(.A(new_n903_), .B(new_n692_), .C1(new_n887_), .C2(new_n889_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n656_), .A2(new_n437_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n270_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n859_), .A2(new_n736_), .A3(new_n389_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G169gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n278_), .A2(new_n279_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n909_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n909_), .A2(G169gat), .A3(new_n911_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n913_), .A2(new_n915_), .A3(new_n916_), .ZN(G1348gat));
  NOR2_X1   g716(.A1(new_n882_), .A2(new_n441_), .ZN(new_n918_));
  AND4_X1   g717(.A1(G176gat), .A2(new_n918_), .A3(new_n587_), .A4(new_n908_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n859_), .A2(new_n908_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n587_), .A3(new_n389_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n921_), .B2(new_n216_), .ZN(G1349gat));
  NOR3_X1   g721(.A1(new_n907_), .A2(new_n640_), .A3(new_n270_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G183gat), .B1(new_n918_), .B2(new_n923_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n920_), .A2(new_n389_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n640_), .A2(new_n231_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n920_), .A2(new_n389_), .A3(new_n622_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G190gat), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n920_), .A2(new_n650_), .A3(new_n232_), .A4(new_n389_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1351gat));
  NOR4_X1   g730(.A1(new_n882_), .A2(new_n439_), .A3(new_n389_), .A4(new_n907_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n736_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT124), .B(G197gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n587_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g736(.A1(new_n883_), .A2(new_n906_), .ZN(new_n938_));
  AND2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n938_), .A2(new_n640_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n932_), .B2(new_n685_), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT125), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n932_), .B(new_n685_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n938_), .A2(new_n640_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n945_), .B(new_n946_), .C1(new_n947_), .C2(new_n940_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n944_), .A2(new_n948_), .ZN(G1354gat));
  NAND3_X1  g748(.A1(new_n883_), .A2(new_n650_), .A3(new_n906_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT126), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n932_), .A2(new_n952_), .A3(new_n650_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n951_), .A2(new_n290_), .A3(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n622_), .A2(G218gat), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n955_), .B(KEYINPUT127), .Z(new_n956_));
  NAND2_X1  g755(.A1(new_n932_), .A2(new_n956_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n954_), .A2(new_n957_), .ZN(G1355gat));
endmodule


