//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n584_, new_n585_, new_n586_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT64), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n217_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n213_), .A2(KEYINPUT64), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT65), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n228_), .B(KEYINPUT7), .Z(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n211_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  AOI211_X1 g030(.A(KEYINPUT66), .B(new_n229_), .C1(new_n220_), .C2(new_n226_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G85gat), .B(G92gat), .Z(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n218_), .B2(new_n219_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n224_), .A2(new_n238_), .A3(new_n225_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n230_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n234_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n233_), .A2(new_n236_), .B1(KEYINPUT8), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G85gat), .ZN(new_n243_));
  INV_X1    g042(.A(G92gat), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT9), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT10), .B(G99gat), .Z(new_n247_));
  INV_X1    g046(.A(G106gat), .ZN(new_n248_));
  AOI22_X1  g047(.A1(KEYINPUT9), .A2(new_n234_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n227_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n208_), .B(new_n210_), .C1(new_n242_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n218_), .A2(new_n219_), .A3(new_n212_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT65), .B1(new_n224_), .B2(new_n225_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n230_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT66), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n227_), .A2(new_n211_), .A3(new_n230_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n236_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n251_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n253_), .B1(new_n261_), .B2(new_n207_), .ZN(new_n262_));
  AND2_X1   g061(.A1(G230gat), .A2(G233gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n261_), .B2(new_n207_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n252_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n252_), .A2(new_n262_), .A3(new_n264_), .A4(KEYINPUT71), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n208_), .B1(new_n242_), .B2(new_n251_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n261_), .A2(new_n271_), .A3(new_n207_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n261_), .B2(new_n207_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n263_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  AND4_X1   g079(.A1(KEYINPUT73), .A2(new_n269_), .A3(new_n275_), .A4(new_n280_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n267_), .A2(new_n268_), .B1(new_n263_), .B2(new_n274_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT73), .B1(new_n282_), .B2(new_n280_), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n281_), .A2(new_n283_), .B1(new_n282_), .B2(new_n280_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT13), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT13), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G29gat), .B(G36gat), .ZN(new_n288_));
  INV_X1    g087(.A(G43gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n288_), .B(G43gat), .ZN(new_n292_));
  INV_X1    g091(.A(G50gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT79), .B(G15gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n297_), .B(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G229gat), .A3(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT15), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n295_), .A2(KEYINPUT74), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n295_), .A2(KEYINPUT74), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT15), .A3(new_n309_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n314_), .A3(new_n305_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n305_), .B2(new_n297_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G229gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT83), .Z(new_n318_));
  OAI21_X1  g117(.A(new_n307_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G113gat), .B(G141gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT85), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G169gat), .ZN(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT84), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n319_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n287_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  OR3_X1    g134(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT94), .ZN(new_n339_));
  INV_X1    g138(.A(G155gat), .ZN(new_n340_));
  INV_X1    g139(.A(G162gat), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT95), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n339_), .B(KEYINPUT1), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(G155gat), .B2(G162gat), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n347_), .B(new_n331_), .C1(G141gat), .C2(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G127gat), .B(G134gat), .ZN(new_n350_));
  INV_X1    g149(.A(G113gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G120gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n349_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n349_), .A2(new_n358_), .A3(new_n353_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n357_), .B1(new_n360_), .B2(new_n356_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT0), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G57gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT105), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n361_), .A2(new_n365_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n361_), .A2(KEYINPUT105), .A3(new_n365_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G204gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(G197gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n323_), .A2(G204gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT21), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n376_), .A2(KEYINPUT99), .A3(G197gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n378_), .A2(KEYINPUT99), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n377_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n379_), .B(new_n380_), .C1(new_n383_), .C2(KEYINPUT21), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT100), .ZN(new_n385_));
  INV_X1    g184(.A(new_n380_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(KEYINPUT21), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT23), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G169gat), .ZN(new_n394_));
  INV_X1    g193(.A(G176gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT87), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G169gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n395_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(KEYINPUT24), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n390_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(KEYINPUT24), .A3(new_n392_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT25), .B(G183gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT26), .B(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n404_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n402_), .A2(new_n405_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n398_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n388_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT20), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n403_), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT104), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n402_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n393_), .A2(new_n396_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n388_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n375_), .B1(new_n413_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n388_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(KEYINPUT20), .C1(new_n411_), .C2(new_n388_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(new_n375_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT18), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G64gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(new_n244_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n423_), .B(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT27), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n427_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n374_), .B1(new_n413_), .B2(new_n419_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n374_), .B2(new_n422_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n434_), .A3(KEYINPUT27), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n437_), .A2(KEYINPUT98), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(KEYINPUT98), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n388_), .A4(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n349_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n443_));
  OAI21_X1  g242(.A(new_n388_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(G228gat), .A3(G233gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G78gat), .B(G106gat), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n447_), .A3(new_n445_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(KEYINPUT102), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n349_), .A2(KEYINPUT29), .A3(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G22gat), .B(G50gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n349_), .B2(KEYINPUT29), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT97), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT97), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n451_), .B(new_n462_), .C1(KEYINPUT102), .C2(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n449_), .A2(new_n458_), .A3(new_n450_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT103), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n449_), .A2(KEYINPUT103), .A3(new_n458_), .A4(new_n450_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n411_), .B(KEYINPUT30), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(G15gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G71gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G99gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT88), .B(G43gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT89), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n476_), .B(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n469_), .A2(new_n470_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT91), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(KEYINPUT92), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n482_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(KEYINPUT92), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n468_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n466_), .A2(new_n467_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n490_), .B1(new_n493_), .B2(new_n463_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n372_), .B(new_n436_), .C1(new_n492_), .C2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n423_), .B1(new_n496_), .B2(new_n428_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n433_), .A2(KEYINPUT32), .A3(new_n427_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n371_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n369_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n369_), .A2(new_n500_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n429_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n356_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n365_), .B1(new_n360_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n504_), .B2(new_n355_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n499_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n468_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n491_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n328_), .B1(new_n495_), .B2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n511_));
  XNOR2_X1  g310(.A(G127gat), .B(G155gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n305_), .B(new_n207_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT81), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT17), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n518_), .A2(new_n515_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n522_), .A2(KEYINPUT17), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n523_), .B2(new_n520_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n312_), .A2(new_n314_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT75), .B1(new_n526_), .B2(new_n261_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n291_), .A2(new_n294_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n261_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n261_), .A2(KEYINPUT75), .A3(new_n528_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n533_), .A2(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G134gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(new_n341_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n544_));
  INV_X1    g343(.A(new_n538_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n530_), .A2(new_n545_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT76), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n546_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n542_), .B(KEYINPUT36), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT77), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT77), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n549_), .A2(new_n553_), .A3(new_n555_), .A4(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT37), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n539_), .A2(KEYINPUT78), .A3(new_n546_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT78), .B1(new_n539_), .B2(new_n546_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n548_), .B1(new_n562_), .B2(new_n551_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n525_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n510_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n300_), .A3(new_n371_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT38), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n563_), .A2(new_n525_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n510_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G1gat), .B1(new_n573_), .B2(new_n372_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(G1324gat));
  INV_X1    g374(.A(new_n436_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n301_), .A3(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G8gat), .B1(new_n573_), .B2(new_n436_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT39), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(KEYINPUT39), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT40), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(G1325gat));
  AOI21_X1  g382(.A(new_n473_), .B1(new_n572_), .B2(new_n490_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT41), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n568_), .A2(new_n473_), .A3(new_n490_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(G1326gat));
  OAI21_X1  g386(.A(G22gat), .B1(new_n573_), .B2(new_n508_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT42), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n508_), .A2(G22gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n567_), .B2(new_n590_), .ZN(G1327gat));
  NAND2_X1  g390(.A1(new_n495_), .A2(new_n509_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n559_), .A2(new_n565_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT43), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n594_), .B2(KEYINPUT106), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n592_), .B(new_n594_), .C1(KEYINPUT106), .C2(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n328_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n525_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT44), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n328_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(KEYINPUT44), .A3(new_n525_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n371_), .A2(G29gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n563_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n524_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n510_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n372_), .ZN(new_n612_));
  OAI22_X1  g411(.A1(new_n607_), .A2(new_n608_), .B1(G29gat), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT107), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1328gat));
  INV_X1    g414(.A(KEYINPUT46), .ZN(new_n616_));
  INV_X1    g415(.A(G36gat), .ZN(new_n617_));
  AND4_X1   g416(.A1(KEYINPUT44), .A2(new_n600_), .A3(new_n601_), .A4(new_n525_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT44), .B1(new_n605_), .B2(new_n525_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n620_), .B2(new_n576_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT45), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n611_), .A2(G36gat), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT108), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n576_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n624_), .B1(new_n623_), .B2(new_n576_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n622_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n627_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(KEYINPUT45), .A3(new_n625_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n616_), .B1(new_n621_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G36gat), .B1(new_n607_), .B2(new_n436_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n633_), .A2(KEYINPUT46), .A3(new_n630_), .A4(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1329gat));
  OAI21_X1  g434(.A(new_n289_), .B1(new_n611_), .B2(new_n491_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT109), .Z(new_n637_));
  NAND2_X1  g436(.A1(new_n490_), .A2(G43gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n607_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g439(.A(new_n293_), .B1(new_n611_), .B2(new_n508_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n468_), .A2(G50gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n607_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT110), .ZN(G1331gat));
  NOR2_X1   g443(.A1(new_n287_), .A2(new_n327_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n592_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n566_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G57gat), .B1(new_n648_), .B2(new_n371_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n571_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT111), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n371_), .A2(G57gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(G1332gat));
  OR3_X1    g453(.A1(new_n647_), .A2(G64gat), .A3(new_n436_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G64gat), .B1(new_n651_), .B2(new_n436_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(G1333gat));
  OR3_X1    g459(.A1(new_n647_), .A2(G71gat), .A3(new_n491_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G71gat), .B1(new_n651_), .B2(new_n491_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT49), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(KEYINPUT49), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(G1334gat));
  OAI21_X1  g464(.A(G78gat), .B1(new_n651_), .B2(new_n508_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT50), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n647_), .A2(G78gat), .A3(new_n508_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1335gat));
  NAND2_X1  g468(.A1(new_n646_), .A2(new_n610_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G85gat), .B1(new_n671_), .B2(new_n371_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n600_), .A2(KEYINPUT113), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n645_), .A2(new_n525_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n600_), .A2(KEYINPUT113), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n673_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n372_), .A2(new_n243_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n672_), .B1(new_n677_), .B2(new_n678_), .ZN(G1336gat));
  AOI21_X1  g478(.A(G92gat), .B1(new_n671_), .B2(new_n576_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n436_), .A2(new_n244_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n677_), .B2(new_n681_), .ZN(G1337gat));
  NAND4_X1  g481(.A1(new_n673_), .A2(new_n490_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G99gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n671_), .A2(new_n247_), .A3(new_n490_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n687_));
  NAND2_X1  g486(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n688_), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1338gat));
  NAND3_X1  g489(.A1(new_n671_), .A2(new_n248_), .A3(new_n468_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n600_), .A2(new_n468_), .A3(new_n675_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT52), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G106gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G106gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g496(.A(new_n280_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n252_), .B(new_n262_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n263_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT55), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n265_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT55), .B1(new_n267_), .B2(new_n268_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT56), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n283_), .B2(new_n281_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n306_), .A2(new_n318_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n708_));
  MUX2_X1   g507(.A(new_n319_), .B(new_n708_), .S(new_n324_), .Z(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n704_), .B2(KEYINPUT56), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n706_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT117), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(KEYINPUT58), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT58), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT117), .B(new_n714_), .C1(new_n706_), .C2(new_n710_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n713_), .A2(new_n565_), .A3(new_n559_), .A4(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT57), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n327_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT115), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n327_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT116), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n704_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n704_), .A2(new_n722_), .A3(KEYINPUT56), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n719_), .A2(new_n721_), .A3(new_n725_), .A4(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n284_), .A2(new_n709_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n717_), .B1(new_n729_), .B2(new_n609_), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT57), .B(new_n563_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n716_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT118), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT118), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n716_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n525_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n327_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n566_), .A2(new_n737_), .A3(new_n287_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT54), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n566_), .A2(new_n740_), .A3(new_n737_), .A4(new_n287_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n736_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n576_), .A2(new_n372_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n492_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT59), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n732_), .A2(new_n525_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n742_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n746_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n748_), .A2(G113gat), .A3(new_n327_), .A4(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT120), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n747_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n745_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT119), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n737_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n760_), .B2(G113gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n758_), .A2(KEYINPUT119), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n758_), .A2(KEYINPUT119), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n327_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(KEYINPUT120), .A3(new_n351_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n754_), .B1(new_n761_), .B2(new_n765_), .ZN(G1340gat));
  INV_X1    g565(.A(new_n287_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n752_), .C1(new_n758_), .C2(new_n751_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT121), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n769_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(G120gat), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n757_), .A2(new_n759_), .ZN(new_n773_));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n773_), .B(new_n775_), .C1(KEYINPUT60), .C2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(G1341gat));
  AOI21_X1  g576(.A(G127gat), .B1(new_n773_), .B2(new_n524_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G127gat), .B1(new_n525_), .B2(KEYINPUT122), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n748_), .B(new_n752_), .C1(KEYINPUT122), .C2(G127gat), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n778_), .B1(new_n779_), .B2(new_n781_), .ZN(G1342gat));
  AOI21_X1  g581(.A(G134gat), .B1(new_n773_), .B2(new_n563_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n748_), .A2(new_n752_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n594_), .A2(G134gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT123), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(G1343gat));
  AND2_X1   g586(.A1(new_n743_), .A2(new_n494_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n744_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n737_), .ZN(new_n790_));
  INV_X1    g589(.A(G141gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1344gat));
  NOR2_X1   g591(.A1(new_n789_), .A2(new_n287_), .ZN(new_n793_));
  INV_X1    g592(.A(G148gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1345gat));
  NOR2_X1   g594(.A1(new_n789_), .A2(new_n525_), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT61), .B(G155gat), .Z(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(G1346gat));
  NOR3_X1   g597(.A1(new_n789_), .A2(new_n341_), .A3(new_n593_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n789_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n563_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n341_), .B2(new_n801_), .ZN(G1347gat));
  INV_X1    g601(.A(KEYINPUT124), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n436_), .A2(new_n371_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n490_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n749_), .B2(new_n742_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n327_), .A3(new_n508_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G169gat), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n806_), .A2(new_n327_), .A3(new_n394_), .A4(new_n508_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT62), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT62), .B1(new_n807_), .B2(G169gat), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n803_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(KEYINPUT124), .A3(new_n812_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1348gat));
  NAND2_X1  g617(.A1(new_n806_), .A2(new_n508_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G176gat), .B1(new_n820_), .B2(new_n767_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n468_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n805_), .A2(new_n395_), .A3(new_n287_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(G1349gat));
  NOR3_X1   g623(.A1(new_n819_), .A2(new_n406_), .A3(new_n525_), .ZN(new_n825_));
  INV_X1    g624(.A(G183gat), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n822_), .A2(new_n490_), .A3(new_n524_), .A4(new_n804_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1350gat));
  NAND3_X1  g627(.A1(new_n820_), .A2(new_n407_), .A3(new_n563_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G190gat), .B1(new_n819_), .B2(new_n593_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1351gat));
  NAND2_X1  g630(.A1(new_n788_), .A2(new_n804_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n737_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(new_n323_), .ZN(G1352gat));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n376_), .A2(KEYINPUT125), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n376_), .A2(KEYINPUT125), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n767_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n832_), .A2(new_n287_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n836_), .ZN(G1353gat));
  NAND3_X1  g639(.A1(new_n788_), .A2(new_n524_), .A3(new_n804_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n842_));
  AND2_X1   g641(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n841_), .B2(new_n842_), .ZN(G1354gat));
  NAND3_X1  g644(.A1(new_n835_), .A2(G218gat), .A3(new_n594_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n743_), .A2(new_n494_), .A3(new_n563_), .A4(new_n804_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n847_), .A2(KEYINPUT126), .ZN(new_n848_));
  INV_X1    g647(.A(G218gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(KEYINPUT126), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n846_), .A2(new_n851_), .ZN(G1355gat));
endmodule


