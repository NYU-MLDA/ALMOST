//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G197gat), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT92), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT21), .B1(new_n204_), .B2(KEYINPUT92), .ZN(new_n209_));
  OAI221_X1 g008(.A(new_n202_), .B1(KEYINPUT21), .B2(new_n207_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(KEYINPUT21), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(new_n202_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G228gat), .A2(G233gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT91), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(KEYINPUT93), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT29), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n219_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n225_), .B(KEYINPUT3), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n227_), .B(KEYINPUT2), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n217_), .B1(new_n218_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n216_), .A2(KEYINPUT93), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI221_X1 g036(.A(new_n217_), .B1(KEYINPUT93), .B2(new_n216_), .C1(new_n218_), .C2(new_n234_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G78gat), .B(G106gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n234_), .B2(new_n218_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G22gat), .B(G50gat), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR4_X1   g044(.A1(new_n229_), .A2(new_n233_), .A3(KEYINPUT29), .A4(new_n241_), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n240_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n239_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AND4_X1   g051(.A1(KEYINPUT94), .A2(new_n237_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(KEYINPUT90), .A3(new_n248_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT90), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n251_), .A2(KEYINPUT94), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n240_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n252_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT19), .ZN(new_n262_));
  NOR2_X1   g061(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G169gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n264_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G183gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT25), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G183gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT26), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT83), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n273_), .A4(new_n275_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n288_), .A2(G169gat), .A3(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT84), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n287_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n270_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT84), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(G169gat), .B2(G176gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n293_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n271_), .B1(new_n286_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT85), .B(new_n271_), .C1(new_n286_), .C2(new_n299_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n213_), .A3(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n210_), .A2(new_n212_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n276_), .A2(new_n281_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n271_), .B1(new_n299_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT95), .B1(new_n304_), .B2(KEYINPUT20), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n262_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n303_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n306_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT20), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n262_), .A2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n314_), .B(new_n316_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT18), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G64gat), .B(G92gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G57gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(new_n233_), .B2(new_n229_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT96), .ZN(new_n334_));
  INV_X1    g133(.A(new_n233_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n330_), .B(new_n331_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n228_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n234_), .A2(KEYINPUT96), .A3(new_n336_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n333_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n329_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n350_), .A2(new_n328_), .A3(new_n347_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n324_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT95), .ZN(new_n354_));
  INV_X1    g153(.A(new_n303_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n296_), .A2(new_n297_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n270_), .B1(new_n287_), .B2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n357_), .A2(new_n282_), .A3(new_n298_), .A4(new_n285_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT85), .B1(new_n358_), .B2(new_n271_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n355_), .A2(new_n359_), .A3(new_n306_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n360_), .B2(new_n315_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n262_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n309_), .A4(new_n305_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT99), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n305_), .A2(new_n309_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n362_), .A4(new_n361_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n306_), .B1(new_n308_), .B2(KEYINPUT98), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(KEYINPUT98), .B2(new_n308_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n314_), .A2(new_n369_), .A3(KEYINPUT20), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n262_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n323_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT100), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(KEYINPUT100), .A3(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n353_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n346_), .A2(new_n329_), .A3(new_n348_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n351_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n343_), .A2(new_n344_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n338_), .A2(new_n339_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n384_), .B(new_n328_), .C1(new_n344_), .C2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n318_), .A2(new_n322_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n312_), .A2(new_n322_), .A3(new_n317_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n260_), .B1(new_n378_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT101), .ZN(new_n393_));
  INV_X1    g192(.A(new_n260_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n349_), .A2(new_n351_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n323_), .B2(new_n318_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n363_), .A2(KEYINPUT99), .B1(new_n262_), .B2(new_n370_), .ZN(new_n397_));
  AOI211_X1 g196(.A(new_n375_), .B(new_n323_), .C1(new_n397_), .C2(new_n367_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT100), .B1(new_n372_), .B2(new_n373_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n396_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n388_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n383_), .A2(new_n386_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n389_), .A4(new_n381_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n394_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT101), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n260_), .A2(new_n352_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n322_), .B1(new_n397_), .B2(new_n367_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n389_), .A2(KEYINPUT27), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT102), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n322_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n372_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT102), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT27), .A4(new_n389_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n407_), .A2(new_n410_), .A3(new_n412_), .A4(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n393_), .A2(new_n406_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT87), .B(G43gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n313_), .B(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT31), .Z(new_n421_));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(G15gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G71gat), .ZN(new_n425_));
  INV_X1    g224(.A(G99gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT86), .B(KEYINPUT30), .Z(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(new_n336_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n421_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT88), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT103), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n410_), .A2(new_n416_), .A3(new_n431_), .A4(new_n412_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n260_), .A2(new_n395_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OR3_X1    g235(.A1(new_n434_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n418_), .A2(new_n432_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G29gat), .B(G36gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n439_), .A2(KEYINPUT71), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(KEYINPUT71), .ZN(new_n441_));
  XOR2_X1   g240(.A(G43gat), .B(G50gat), .Z(new_n442_));
  OR3_X1    g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G15gat), .B(G22gat), .ZN(new_n448_));
  INV_X1    g247(.A(G1gat), .ZN(new_n449_));
  INV_X1    g248(.A(G8gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT14), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G1gat), .B(G8gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n447_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n445_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n464_), .A2(KEYINPUT81), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n459_), .B(new_n445_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n464_), .B(KEYINPUT81), .C1(new_n463_), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G113gat), .B(G141gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G169gat), .B(G197gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n465_), .A2(new_n467_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(KEYINPUT82), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n438_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT104), .ZN(new_n482_));
  OR3_X1    g281(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT7), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT6), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(KEYINPUT7), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT10), .B(G99gat), .Z(new_n493_));
  INV_X1    g292(.A(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n496_));
  INV_X1    g295(.A(G85gat), .ZN(new_n497_));
  INV_X1    g296(.A(G92gat), .ZN(new_n498_));
  OR3_X1    g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT9), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n496_), .A3(new_n486_), .A4(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT65), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n492_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n447_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n491_), .A2(new_n492_), .A3(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n445_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT73), .B1(new_n502_), .B2(new_n447_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n508_), .A2(KEYINPUT35), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n508_), .A2(KEYINPUT35), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n503_), .B(new_n505_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n505_), .A2(new_n503_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n519_), .B(KEYINPUT36), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n521_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT37), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n516_), .B2(KEYINPUT74), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n513_), .A2(new_n527_), .A3(new_n515_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n526_), .A2(new_n528_), .B1(new_n520_), .B2(new_n516_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n529_), .A2(KEYINPUT75), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT75), .B1(new_n529_), .B2(new_n530_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n525_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n537_));
  XOR2_X1   g336(.A(G71gat), .B(G78gat), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n504_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(KEYINPUT67), .Z(new_n543_));
  NAND3_X1  g342(.A1(new_n502_), .A2(new_n543_), .A3(KEYINPUT12), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n541_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT12), .B1(new_n502_), .B2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT64), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n502_), .A2(new_n546_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n542_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G176gat), .B(G204gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT69), .ZN(new_n557_));
  XOR2_X1   g356(.A(G120gat), .B(G148gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(KEYINPUT70), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n555_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n459_), .B(new_n570_), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT80), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(new_n541_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n541_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT17), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(KEYINPUT17), .ZN(new_n581_));
  OR4_X1    g380(.A1(new_n573_), .A2(new_n574_), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n571_), .A2(new_n543_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n571_), .A2(new_n543_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT79), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(KEYINPUT79), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n582_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n534_), .A2(new_n569_), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n482_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n449_), .A3(new_n352_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n569_), .A2(new_n588_), .A3(new_n529_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n481_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n395_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n592_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n597_), .A3(new_n598_), .ZN(G1324gat));
  AND3_X1   g398(.A1(new_n416_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n590_), .A2(new_n450_), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT105), .B1(new_n596_), .B2(new_n600_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT105), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n604_), .A3(new_n601_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(G8gat), .A3(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT39), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT39), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n602_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT40), .B(new_n602_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1325gat));
  INV_X1    g412(.A(new_n432_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n423_), .B1(new_n595_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n590_), .A2(new_n423_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n595_), .B2(new_n394_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n590_), .A2(new_n619_), .A3(new_n394_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n569_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n588_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n529_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n482_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n352_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n588_), .A3(new_n479_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n417_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT101), .B(new_n394_), .C1(new_n400_), .C2(new_n403_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n432_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n437_), .A2(new_n436_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n632_), .B1(new_n637_), .B2(new_n534_), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT43), .B(new_n533_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT44), .B(new_n631_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT43), .B1(new_n438_), .B2(new_n533_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(new_n534_), .A3(new_n632_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n630_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n645_), .B2(KEYINPUT44), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n631_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT106), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n641_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n352_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n629_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  INV_X1    g451(.A(KEYINPUT46), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n650_), .A2(new_n601_), .ZN(new_n654_));
  INV_X1    g453(.A(G36gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n482_), .A2(new_n655_), .A3(new_n601_), .A4(new_n627_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n653_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n657_), .B(new_n658_), .Z(new_n661_));
  OAI211_X1 g460(.A(new_n661_), .B(KEYINPUT46), .C1(new_n654_), .C2(new_n655_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1329gat));
  AND2_X1   g462(.A1(new_n431_), .A2(G43gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n650_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n650_), .A2(KEYINPUT108), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n628_), .A2(new_n614_), .ZN(new_n669_));
  INV_X1    g468(.A(G43gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT47), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n667_), .A2(new_n674_), .A3(new_n668_), .A4(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1330gat));
  INV_X1    g475(.A(G50gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n628_), .A2(new_n677_), .A3(new_n394_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n640_), .A2(new_n394_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n645_), .A2(new_n642_), .A3(KEYINPUT44), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT106), .B1(new_n647_), .B2(new_n648_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n679_), .B1(new_n684_), .B2(G50gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n680_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(KEYINPUT109), .A3(new_n677_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n678_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT110), .B(new_n678_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1331gat));
  INV_X1    g491(.A(G57gat), .ZN(new_n693_));
  INV_X1    g492(.A(new_n588_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n637_), .A2(new_n569_), .A3(new_n694_), .A4(new_n480_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n533_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n697_), .B2(new_n395_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT111), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n626_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n700_), .A2(new_n693_), .A3(new_n395_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n700_), .B2(new_n600_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n600_), .A2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n697_), .B2(new_n705_), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n700_), .B2(new_n432_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT49), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n432_), .A2(G71gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n697_), .B2(new_n709_), .ZN(G1334gat));
  OR3_X1    g509(.A1(new_n697_), .A2(G78gat), .A3(new_n260_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G78gat), .B1(new_n700_), .B2(new_n260_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT113), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n713_), .A2(new_n715_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n711_), .B1(new_n716_), .B2(new_n717_), .ZN(G1335gat));
  NAND2_X1  g517(.A1(new_n569_), .A2(new_n588_), .ZN(new_n719_));
  NOR4_X1   g518(.A1(new_n438_), .A2(new_n719_), .A3(new_n626_), .A4(new_n479_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n497_), .A3(new_n352_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n479_), .B(new_n719_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n352_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n497_), .ZN(G1336gat));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n498_), .A3(new_n601_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n722_), .A2(new_n601_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n498_), .ZN(G1337gat));
  NAND3_X1  g526(.A1(new_n720_), .A2(new_n493_), .A3(new_n431_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT114), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n426_), .B1(new_n722_), .B2(new_n614_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g531(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n722_), .A2(new_n394_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G106gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT52), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n720_), .A2(new_n494_), .A3(new_n394_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(KEYINPUT52), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n734_), .B2(G106gat), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n737_), .B(new_n733_), .C1(new_n739_), .C2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n738_), .A2(new_n743_), .ZN(G1339gat));
  XNOR2_X1  g543(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n589_), .B2(new_n480_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n589_), .A2(new_n480_), .ZN(new_n747_));
  AND2_X1   g546(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n551_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT55), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n551_), .A2(new_n750_), .A3(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n752_), .B(new_n754_), .C1(new_n550_), .C2(new_n548_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n563_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT56), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n758_), .A3(new_n563_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n757_), .A2(new_n479_), .A3(new_n562_), .A4(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n466_), .B1(G229gat), .B2(G233gat), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n761_), .A2(KEYINPUT118), .A3(new_n471_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT118), .B1(new_n761_), .B2(new_n471_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n462_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n762_), .B(new_n763_), .C1(new_n463_), .C2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n472_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n565_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n529_), .B1(new_n760_), .B2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT57), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n757_), .A2(new_n562_), .A3(new_n766_), .A4(new_n759_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT58), .B1(new_n770_), .B2(KEYINPUT119), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n756_), .A2(KEYINPUT56), .B1(new_n555_), .B2(new_n561_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n766_), .A4(new_n759_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n533_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n772_), .B1(new_n777_), .B2(KEYINPUT120), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n770_), .A2(KEYINPUT119), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n771_), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n534_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n769_), .B1(new_n778_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n749_), .B1(new_n784_), .B2(new_n694_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n434_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n479_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(KEYINPUT59), .A3(new_n786_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n480_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n794_), .B2(new_n789_), .ZN(G1340gat));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n624_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n788_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n796_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n624_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n796_), .ZN(G1341gat));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n788_), .A2(new_n801_), .A3(new_n694_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n588_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n801_), .ZN(G1342gat));
  AOI21_X1  g603(.A(G134gat), .B1(new_n788_), .B2(new_n529_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n792_), .A2(new_n793_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n534_), .A2(G134gat), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT121), .Z(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n806_), .B2(new_n808_), .ZN(G1343gat));
  NOR3_X1   g608(.A1(new_n614_), .A2(new_n260_), .A3(new_n395_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n785_), .A2(new_n600_), .A3(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n480_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n624_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g614(.A1(new_n811_), .A2(new_n588_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT61), .B(G155gat), .Z(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1346gat));
  INV_X1    g617(.A(G162gat), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n811_), .A2(new_n819_), .A3(new_n533_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n811_), .B2(new_n626_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT122), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(new_n819_), .C1(new_n811_), .C2(new_n626_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n820_), .B1(new_n822_), .B2(new_n824_), .ZN(G1347gat));
  NOR2_X1   g624(.A1(new_n432_), .A2(new_n435_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n785_), .A2(new_n479_), .A3(new_n601_), .A4(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT62), .B1(new_n827_), .B2(KEYINPUT22), .ZN(new_n828_));
  OAI21_X1  g627(.A(G169gat), .B1(new_n827_), .B2(KEYINPUT62), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n290_), .B2(new_n828_), .ZN(G1348gat));
  NAND2_X1  g630(.A1(KEYINPUT123), .A2(G176gat), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n785_), .A2(new_n601_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n826_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n834_), .B2(new_n624_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT123), .B(G176gat), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n833_), .A2(new_n569_), .A3(new_n826_), .A4(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1349gat));
  OAI21_X1  g637(.A(new_n272_), .B1(new_n834_), .B2(new_n588_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n833_), .A2(new_n694_), .A3(new_n276_), .A4(new_n826_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1350gat));
  OAI21_X1  g640(.A(G190gat), .B1(new_n834_), .B2(new_n533_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n529_), .A2(new_n283_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n834_), .B2(new_n843_), .ZN(G1351gat));
  AND2_X1   g643(.A1(new_n432_), .A2(new_n407_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n833_), .A2(new_n479_), .A3(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g646(.A1(new_n785_), .A2(new_n569_), .A3(new_n601_), .A4(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT125), .B1(new_n849_), .B2(G204gat), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n848_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT126), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT126), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n852_), .B(new_n857_), .C1(new_n848_), .C2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1353gat));
  NAND3_X1  g658(.A1(new_n833_), .A2(new_n694_), .A3(new_n845_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT63), .B(G211gat), .Z(new_n863_));
  NAND4_X1  g662(.A1(new_n833_), .A2(new_n694_), .A3(new_n845_), .A4(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1354gat));
  AND2_X1   g664(.A1(new_n833_), .A2(new_n845_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT127), .B(G218gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n533_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n833_), .A2(new_n529_), .A3(new_n845_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n866_), .A2(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1355gat));
endmodule


