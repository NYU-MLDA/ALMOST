//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  OAI211_X1 g009(.A(G85gat), .B(G92gat), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n211_));
  OAI211_X1 g010(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n211_), .B(new_n212_), .Z(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(G106gat), .ZN(new_n215_));
  OR3_X1    g014(.A1(new_n213_), .A2(new_n208_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G29gat), .B(G36gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT68), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n219_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n221_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G232gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT34), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT67), .B(KEYINPUT35), .Z(new_n232_));
  AOI22_X1  g031(.A1(new_n218_), .A2(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n222_), .A2(new_n226_), .A3(KEYINPUT15), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT15), .B1(new_n222_), .B2(new_n226_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n217_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(new_n232_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n233_), .B(new_n236_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G190gat), .B(G218gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G134gat), .B(G162gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT36), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n247_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n241_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n248_), .B(KEYINPUT71), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n239_), .A3(new_n240_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT84), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT21), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(G197gat), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n264_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n268_), .B1(new_n276_), .B2(G197gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT83), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n263_), .B1(new_n272_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G197gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n280_), .A3(new_n264_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(G197gat), .B2(G204gat), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n282_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n261_), .B1(new_n277_), .B2(KEYINPUT21), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT82), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n265_), .A2(new_n266_), .A3(G197gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n284_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT81), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n262_), .B1(new_n270_), .B2(new_n283_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n279_), .B1(new_n289_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(KEYINPUT1), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306_));
  INV_X1    g105(.A(new_n303_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n305_), .A2(KEYINPUT77), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n303_), .C1(new_n304_), .C2(KEYINPUT1), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n302_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n303_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n301_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n299_), .B2(KEYINPUT78), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n299_), .A2(KEYINPUT78), .A3(new_n318_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n313_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n311_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT79), .B1(new_n298_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n279_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n294_), .A2(new_n296_), .A3(new_n295_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n296_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331_));
  INV_X1    g130(.A(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT29), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n326_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n326_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n260_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n323_), .A2(new_n324_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT28), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  NOR2_X1   g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n326_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n338_), .B1(new_n326_), .B2(new_n334_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT85), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n337_), .A2(new_n349_), .A3(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n350_), .A3(new_n258_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353_));
  INV_X1    g152(.A(G43gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(G15gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n355_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT23), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(G183gat), .B2(G190gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G190gat), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n366_), .A2(KEYINPUT75), .A3(KEYINPUT26), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT26), .B1(new_n366_), .B2(KEYINPUT75), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G169gat), .ZN(new_n373_));
  INV_X1    g172(.A(G176gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OR3_X1    g174(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n370_), .A2(new_n361_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n365_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT30), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n379_), .A2(KEYINPUT76), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(KEYINPUT76), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n359_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n359_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G127gat), .B(G134gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G120gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n387_), .B(KEYINPUT31), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n384_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n384_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n382_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT87), .ZN(new_n394_));
  INV_X1    g193(.A(new_n387_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n311_), .B2(new_n322_), .ZN(new_n396_));
  INV_X1    g195(.A(G141gat), .ZN(new_n397_));
  INV_X1    g196(.A(G148gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT78), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT3), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(new_n321_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n303_), .A3(new_n312_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n305_), .A2(KEYINPUT77), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n307_), .A2(new_n306_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n403_), .A2(new_n310_), .A3(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n402_), .B(new_n387_), .C1(new_n405_), .C2(new_n302_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n394_), .B1(new_n396_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n396_), .A2(new_n406_), .A3(KEYINPUT4), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n395_), .B(new_n410_), .C1(new_n311_), .C2(new_n322_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n394_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n408_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT88), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT0), .B(G57gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n414_), .A2(KEYINPUT95), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n413_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n421_), .A2(new_n419_), .A3(new_n407_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n421_), .B2(new_n407_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT95), .A3(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n389_), .A2(new_n392_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n337_), .A2(new_n260_), .A3(new_n339_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n344_), .B1(new_n427_), .B2(new_n340_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n352_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT19), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n378_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT20), .B1(new_n298_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n368_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(new_n375_), .A3(new_n361_), .A4(new_n376_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n365_), .A2(new_n438_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n279_), .B(new_n439_), .C1(new_n289_), .C2(new_n297_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n433_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n330_), .A2(new_n439_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n327_), .B(new_n434_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(KEYINPUT20), .A3(new_n432_), .A4(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT18), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n444_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(KEYINPUT86), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453_));
  AOI211_X1 g252(.A(new_n453_), .B(new_n449_), .C1(new_n441_), .C2(new_n444_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n430_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n451_), .A2(new_n430_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n442_), .A2(KEYINPUT20), .A3(new_n443_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(new_n432_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n439_), .B(KEYINPUT93), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT20), .B1(new_n459_), .B2(new_n330_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT94), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n330_), .A2(new_n378_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT94), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(KEYINPUT20), .C1(new_n459_), .C2(new_n330_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n465_), .B2(new_n432_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n456_), .B1(new_n466_), .B2(new_n448_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n455_), .A2(KEYINPUT96), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT96), .B1(new_n455_), .B2(new_n467_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n429_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT97), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT97), .B(new_n429_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n389_), .A2(new_n392_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n352_), .A2(new_n428_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n448_), .A2(KEYINPUT32), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n465_), .A2(new_n432_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n458_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n441_), .A2(new_n444_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n478_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n420_), .A2(new_n483_), .A3(new_n424_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n452_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n423_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT90), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n423_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n409_), .A2(new_n413_), .A3(new_n411_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT91), .ZN(new_n493_));
  INV_X1    g292(.A(new_n396_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n406_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n419_), .B1(new_n496_), .B2(new_n394_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n489_), .A2(new_n491_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n451_), .A2(KEYINPUT86), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n414_), .A2(KEYINPUT89), .A3(KEYINPUT33), .A4(new_n419_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n501_), .B1(new_n423_), .B2(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n486_), .A2(new_n498_), .A3(new_n499_), .A4(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n485_), .B1(new_n504_), .B2(KEYINPUT92), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n493_), .A2(new_n497_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n423_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n490_), .B1(new_n423_), .B2(new_n487_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n500_), .A2(new_n502_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n452_), .A2(new_n454_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n477_), .B1(new_n505_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n420_), .A2(new_n424_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n477_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n455_), .A2(new_n467_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n476_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n520_));
  AOI211_X1 g319(.A(KEYINPUT99), .B(new_n257_), .C1(new_n474_), .C2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT99), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n455_), .A2(KEYINPUT96), .A3(new_n467_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT97), .B1(new_n526_), .B2(new_n429_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n473_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n482_), .A2(new_n448_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n453_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(new_n499_), .A3(new_n450_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n503_), .B(new_n506_), .C1(new_n508_), .C2(new_n507_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT92), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n481_), .A2(new_n484_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n514_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n340_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n426_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n537_), .A2(new_n344_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n516_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n518_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n535_), .A2(new_n538_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n527_), .A2(new_n528_), .B1(new_n542_), .B2(new_n475_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n522_), .B1(new_n543_), .B2(new_n256_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n521_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT11), .Z(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT65), .B(G71gat), .ZN(new_n548_));
  INV_X1    g347(.A(G78gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(KEYINPUT11), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n217_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n210_), .A2(new_n216_), .A3(new_n551_), .A4(new_n553_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT12), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n217_), .A2(new_n558_), .A3(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G120gat), .B(G148gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n562_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n561_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n573_), .B2(new_n563_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT13), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT74), .ZN(new_n579_));
  INV_X1    g378(.A(G22gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n357_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G15gat), .A2(G22gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G1gat), .A2(G8gat), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n581_), .A2(new_n582_), .B1(KEYINPUT14), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n579_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n227_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n579_), .B(new_n584_), .Z(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n590_), .B2(new_n228_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n234_), .A2(new_n235_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n589_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n590_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n554_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n604_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n604_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n577_), .A2(new_n601_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n545_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n539_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G1gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n601_), .B1(new_n474_), .B2(new_n520_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n250_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n256_), .A2(new_n620_), .A3(KEYINPUT37), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n250_), .B(new_n255_), .C1(new_n619_), .C2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n613_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n577_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n618_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n618_), .A2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT98), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n516_), .A2(G1gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n617_), .A2(new_n636_), .A3(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  INV_X1    g438(.A(new_n526_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(new_n614_), .C1(new_n521_), .C2(new_n544_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n642_), .A3(G8gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n641_), .B2(G8gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n639_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(G8gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT101), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n642_), .A3(G8gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT39), .A3(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n526_), .A2(G8gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n630_), .A2(new_n632_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n630_), .A2(KEYINPUT100), .A3(new_n632_), .A4(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n645_), .A2(new_n649_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n645_), .A2(new_n649_), .A3(KEYINPUT40), .A4(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  NAND3_X1  g459(.A1(new_n628_), .A2(new_n357_), .A3(new_n475_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n545_), .A2(new_n475_), .A3(new_n614_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT41), .B1(new_n662_), .B2(G15gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT102), .B(new_n661_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n538_), .B(KEYINPUT103), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n615_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n672_), .B2(G22gat), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT42), .B(new_n580_), .C1(new_n615_), .C2(new_n671_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n580_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT104), .Z(new_n676_));
  OAI22_X1  g475(.A1(new_n673_), .A2(new_n674_), .B1(new_n631_), .B2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(new_n624_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n543_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n625_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n577_), .A2(new_n601_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n543_), .A2(KEYINPUT43), .A3(new_n678_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n682_), .A4(new_n683_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n539_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G29gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n625_), .A2(new_n256_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n577_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n618_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n516_), .A2(G29gat), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT105), .Z(new_n696_));
  OAI21_X1  g495(.A(new_n690_), .B1(new_n694_), .B2(new_n696_), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n686_), .A2(new_n640_), .A3(new_n687_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G36gat), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n694_), .A2(G36gat), .A3(new_n526_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT45), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(new_n701_), .A3(KEYINPUT46), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n686_), .A2(G43gat), .A3(new_n475_), .A4(new_n687_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n354_), .B1(new_n694_), .B2(new_n476_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g509(.A(G50gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n538_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n618_), .A2(new_n671_), .A3(new_n693_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n688_), .A2(new_n712_), .B1(new_n711_), .B2(new_n713_), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n543_), .A2(new_n601_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT106), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n543_), .A2(new_n717_), .A3(new_n601_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n577_), .A3(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n626_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n539_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n599_), .A2(new_n600_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n576_), .A2(new_n722_), .A3(new_n613_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(G57gat), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n545_), .A2(new_n539_), .A3(new_n723_), .A4(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n726_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n526_), .A2(G64gat), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n720_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n545_), .A2(new_n640_), .A3(new_n723_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(G64gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n733_), .B2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT110), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n739_), .B(new_n732_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1333gat));
  NOR2_X1   g540(.A1(new_n476_), .A2(G71gat), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n720_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n545_), .A2(new_n475_), .A3(new_n723_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(G71gat), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G71gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT113), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n744_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n720_), .A2(new_n549_), .A3(new_n671_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n545_), .A2(new_n671_), .A3(new_n723_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(G78gat), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT115), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n719_), .A2(new_n692_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n539_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n679_), .A2(new_n680_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n576_), .A2(new_n722_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(new_n613_), .A3(new_n683_), .A4(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT116), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n681_), .A2(new_n770_), .A3(new_n683_), .A4(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n539_), .A2(G85gat), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT117), .Z(new_n774_));
  AOI21_X1  g573(.A(new_n765_), .B1(new_n772_), .B2(new_n774_), .ZN(G1336gat));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n764_), .A2(new_n776_), .A3(new_n640_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n526_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n776_), .ZN(G1337gat));
  NOR2_X1   g578(.A1(new_n476_), .A2(new_n214_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n764_), .A2(new_n780_), .B1(new_n781_), .B2(KEYINPUT51), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n476_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n783_));
  INV_X1    g582(.A(G99gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n781_), .A2(KEYINPUT51), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n785_), .B(new_n787_), .ZN(G1338gat));
  INV_X1    g587(.A(G106gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n764_), .A2(new_n789_), .A3(new_n477_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n681_), .A2(new_n477_), .A3(new_n683_), .A4(new_n767_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(G106gat), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n791_), .B2(G106gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n790_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g596(.A1(new_n640_), .A2(new_n516_), .A3(new_n476_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n573_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n601_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n571_), .A2(new_n722_), .A3(KEYINPUT119), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n557_), .A2(new_n572_), .A3(new_n559_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n562_), .A2(KEYINPUT55), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n570_), .B1(new_n573_), .B2(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n806_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n801_), .B(new_n802_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n600_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n587_), .B1(new_n590_), .B2(new_n228_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n592_), .B2(new_n590_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n597_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n575_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n817_), .A2(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n256_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n816_), .A2(new_n820_), .B1(new_n817_), .B2(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(KEYINPUT57), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n819_), .C1(new_n809_), .C2(new_n815_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n814_), .A2(new_n571_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n828_), .B2(new_n808_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n827_), .B(KEYINPUT56), .C1(new_n804_), .C2(new_n806_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT58), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n804_), .A2(new_n806_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n827_), .A3(new_n826_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n830_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .A4(new_n825_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n678_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n625_), .B1(new_n824_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n624_), .A2(new_n576_), .A3(new_n601_), .A4(new_n625_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n538_), .B(new_n798_), .C1(new_n841_), .C2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n722_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(KEYINPUT122), .A3(new_n849_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n571_), .A2(new_n722_), .A3(KEYINPUT119), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT119), .B1(new_n571_), .B2(new_n722_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n834_), .A2(new_n826_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n853_), .A2(new_n854_), .B1(new_n575_), .B2(new_n814_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n822_), .B1(new_n855_), .B2(new_n819_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n816_), .A2(new_n817_), .A3(KEYINPUT57), .A4(new_n256_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n624_), .B1(new_n831_), .B2(new_n838_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n613_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n842_), .B(KEYINPUT54), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n477_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n798_), .A4(new_n864_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n850_), .A2(new_n865_), .A3(KEYINPUT123), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT123), .B1(new_n850_), .B2(new_n865_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n601_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n848_), .B1(new_n870_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n576_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n846_), .B(new_n873_), .C1(KEYINPUT60), .C2(new_n872_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n576_), .B1(new_n850_), .B2(new_n865_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n872_), .ZN(G1341gat));
  INV_X1    g675(.A(G127gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n846_), .A2(new_n877_), .A3(new_n625_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n613_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n877_), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n624_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n845_), .B2(new_n256_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(KEYINPUT124), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT124), .B1(new_n883_), .B2(new_n884_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1343gat));
  AOI21_X1  g686(.A(new_n475_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n888_));
  AND4_X1   g687(.A1(new_n539_), .A2(new_n888_), .A3(new_n477_), .A4(new_n526_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n722_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n577_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n625_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n889_), .A2(new_n897_), .A3(new_n257_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n889_), .A2(new_n678_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1347gat));
  NAND2_X1  g699(.A1(new_n640_), .A2(new_n425_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n671_), .B(new_n901_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n722_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n373_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(KEYINPUT125), .A3(new_n722_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT22), .B(G169gat), .Z(new_n910_));
  OAI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n903_), .B2(new_n910_), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n902_), .B2(new_n577_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n477_), .B(new_n901_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n576_), .A2(new_n374_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  AOI21_X1  g714(.A(G183gat), .B1(new_n913_), .B2(new_n625_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n613_), .A2(new_n368_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n902_), .B2(new_n917_), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n902_), .A2(new_n436_), .A3(new_n257_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n902_), .A2(new_n678_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n366_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n526_), .A2(new_n517_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n888_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n601_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n280_), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n576_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(G204gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n276_), .B2(new_n926_), .ZN(G1353gat));
  NOR2_X1   g727(.A1(new_n923_), .A2(new_n613_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  AND2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(new_n929_), .B2(new_n930_), .ZN(G1354gat));
  NOR3_X1   g732(.A1(new_n923_), .A2(G218gat), .A3(new_n256_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n923_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n678_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(G218gat), .B2(new_n936_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


