//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_, new_n991_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT8), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT64), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n208_), .B(new_n210_), .C1(new_n215_), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n212_), .A2(new_n214_), .ZN(new_n223_));
  OR2_X1    g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n218_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n205_), .A2(KEYINPUT9), .A3(new_n206_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n219_), .A2(new_n220_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n207_), .B1(new_n230_), .B2(new_n223_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT64), .B(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n222_), .B(new_n229_), .C1(new_n231_), .C2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G78gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT11), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(KEYINPUT11), .B2(new_n235_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n244_), .B2(new_n239_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n208_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n232_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n245_), .A2(new_n247_), .A3(new_n222_), .A4(new_n229_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G230gat), .A2(G233gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n234_), .A2(new_n242_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT12), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT65), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254_));
  AOI211_X1 g053(.A(new_n254_), .B(KEYINPUT12), .C1(new_n234_), .C2(new_n242_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n249_), .B(new_n250_), .C1(new_n253_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n248_), .A2(new_n251_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G230gat), .A3(G233gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G120gat), .B(G148gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT5), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G176gat), .B(G204gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n259_), .B(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT66), .ZN(new_n265_));
  INV_X1    g064(.A(new_n263_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n259_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n202_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G15gat), .ZN(new_n274_));
  INV_X1    g073(.A(G22gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G15gat), .A2(G22gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G1gat), .A2(G8gat), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n276_), .A2(new_n277_), .B1(KEYINPUT14), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n273_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G36gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G29gat), .ZN(new_n282_));
  INV_X1    g081(.A(G29gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G36gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G50gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G43gat), .ZN(new_n287_));
  INV_X1    g086(.A(G43gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G50gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n282_), .A2(new_n284_), .A3(new_n287_), .A4(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n280_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT15), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT15), .B1(new_n291_), .B2(new_n292_), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n280_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n280_), .A2(new_n293_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n295_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G141gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G169gat), .B(G197gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT74), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n303_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n267_), .A2(new_n268_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n264_), .A2(KEYINPUT66), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT13), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n270_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT2), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT3), .B1(new_n319_), .B2(KEYINPUT83), .ZN(new_n320_));
  OR2_X1    g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT82), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n317_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n316_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(KEYINPUT1), .B2(new_n325_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G127gat), .B(G134gat), .Z(new_n336_));
  INV_X1    g135(.A(G120gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G113gat), .ZN(new_n338_));
  INV_X1    g137(.A(G113gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G120gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(KEYINPUT79), .A3(new_n344_), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n336_), .A2(new_n341_), .A3(KEYINPUT79), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n335_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n333_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n342_), .A2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n315_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT4), .B1(new_n335_), .B2(new_n347_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n351_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(KEYINPUT4), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n355_), .B2(new_n315_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n329_), .A2(new_n334_), .A3(new_n350_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n329_), .A2(new_n334_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT4), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n348_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n315_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n352_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n361_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT94), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G183gat), .ZN(new_n379_));
  INV_X1    g178(.A(G190gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT23), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(G183gat), .A3(G190gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT24), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n381_), .A2(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n388_), .A2(KEYINPUT24), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT25), .B(G183gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n386_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n383_), .A2(KEYINPUT77), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n399_), .A2(new_n382_), .A3(G183gat), .A4(G190gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n381_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  INV_X1    g203(.A(G176gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n390_), .B(KEYINPUT95), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n395_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G204gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT87), .B1(new_n411_), .B2(G197gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413_));
  INV_X1    g212(.A(G197gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(G204gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT21), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(G197gat), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n412_), .A2(new_n415_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n411_), .A2(G197gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n414_), .A2(G204gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT21), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G218gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G211gat), .ZN(new_n423_));
  INV_X1    g222(.A(G211gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G218gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n418_), .B(new_n421_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n425_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT88), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n412_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n432_), .A2(KEYINPUT21), .A3(new_n433_), .A4(new_n427_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n410_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n381_), .A2(new_n383_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n397_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G169gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT25), .B1(new_n379_), .B2(KEYINPUT75), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n379_), .A2(KEYINPUT25), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n392_), .B(new_n443_), .C1(new_n444_), .C2(KEYINPUT75), .ZN(new_n445_));
  INV_X1    g244(.A(new_n389_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(KEYINPUT76), .A2(G169gat), .A3(G176gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n384_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n448_), .A3(new_n391_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n402_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n442_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n435_), .A2(KEYINPUT89), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n430_), .A2(new_n434_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n451_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n378_), .B1(new_n437_), .B2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G8gat), .B(G36gat), .Z(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n410_), .B2(new_n436_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n452_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n377_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(new_n461_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT101), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT101), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n456_), .A2(new_n465_), .A3(new_n468_), .A4(new_n461_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n461_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n437_), .A2(new_n455_), .A3(new_n378_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n377_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n467_), .A2(KEYINPUT27), .A3(new_n469_), .A4(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n463_), .A2(new_n377_), .A3(new_n464_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n451_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n454_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n453_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n386_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n450_), .A2(new_n396_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n408_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n462_), .B1(new_n482_), .B2(new_n435_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n377_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n470_), .B1(new_n475_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n466_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT27), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n373_), .A2(new_n474_), .A3(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT92), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493_));
  INV_X1    g292(.A(new_n328_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n321_), .B2(new_n318_), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n496_), .A2(KEYINPUT3), .B1(new_n321_), .B2(new_n322_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n497_), .B2(new_n317_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n493_), .B(KEYINPUT29), .C1(new_n498_), .C2(new_n333_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT90), .B1(new_n349_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n501_), .A3(new_n435_), .ZN(new_n502_));
  INV_X1    g301(.A(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(G228gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(G228gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(KEYINPUT91), .A3(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n508_), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n492_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n502_), .A2(KEYINPUT91), .A3(new_n508_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT91), .B1(new_n502_), .B2(new_n508_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n492_), .B(new_n515_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G22gat), .B(G50gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n349_), .A2(new_n524_), .A3(new_n500_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n349_), .B2(new_n500_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n523_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n523_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n522_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n528_), .A2(new_n531_), .A3(new_n522_), .ZN(new_n533_));
  OAI22_X1  g332(.A1(new_n516_), .A2(new_n520_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n491_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(new_n532_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n519_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n451_), .A2(KEYINPUT30), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n442_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G15gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n545_), .B(new_n274_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n288_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G71gat), .B(G99gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n552_), .A2(KEYINPUT78), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n540_), .B1(new_n544_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT78), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n551_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT78), .B1(new_n552_), .B2(new_n553_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n541_), .A4(new_n543_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n347_), .B(KEYINPUT31), .Z(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n489_), .B1(new_n539_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n564_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT81), .A3(new_n562_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n534_), .A2(new_n538_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT97), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT33), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n360_), .B(new_n576_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n348_), .A2(new_n351_), .A3(new_n315_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n360_), .B(new_n579_), .C1(new_n355_), .C2(new_n315_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n485_), .A2(new_n580_), .A3(new_n466_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT98), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n576_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n369_), .A2(new_n370_), .A3(new_n574_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n485_), .A2(new_n466_), .A3(new_n580_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n461_), .A2(KEYINPUT32), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n456_), .A2(new_n465_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT99), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n456_), .A2(new_n465_), .A3(new_n592_), .A4(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n589_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT100), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n598_), .B(new_n595_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n594_), .A2(new_n372_), .A3(new_n597_), .A4(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n582_), .A2(new_n588_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n571_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n566_), .A2(new_n572_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n313_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT35), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT34), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT67), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT67), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT34), .ZN(new_n613_));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n611_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n609_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT69), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT69), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n619_), .B(new_n609_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n615_), .A2(new_n616_), .A3(new_n609_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n618_), .A2(new_n620_), .B1(KEYINPUT70), .B2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n247_), .A2(new_n293_), .A3(new_n222_), .A4(new_n229_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n298_), .A2(new_n299_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT68), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n234_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n234_), .B2(new_n625_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT70), .ZN(new_n631_));
  INV_X1    g430(.A(new_n621_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n631_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n624_), .B(new_n634_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n635_));
  AOI211_X1 g434(.A(KEYINPUT36), .B(new_n608_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n608_), .B(KEYINPUT36), .Z(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n635_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n234_), .A2(new_n625_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT68), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n627_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n634_), .B1(new_n643_), .B2(new_n624_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT71), .B1(new_n640_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT71), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n633_), .A2(new_n646_), .A3(new_n635_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n639_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT72), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n637_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT72), .B(new_n639_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n605_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n633_), .A2(new_n638_), .A3(new_n635_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n637_), .A2(KEYINPUT37), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n245_), .B(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(new_n280_), .ZN(new_n658_));
  XOR2_X1   g457(.A(G127gat), .B(G155gat), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT16), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G183gat), .B(G211gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT17), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n662_), .B(new_n663_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n658_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n655_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n604_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G1gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n372_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT38), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n313_), .A2(new_n669_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n650_), .A2(new_n651_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n603_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT102), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n373_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n674_), .B1(new_n683_), .B2(new_n672_), .ZN(G1324gat));
  INV_X1    g483(.A(G8gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n474_), .A2(new_n488_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n671_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n679_), .A2(new_n686_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G8gat), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT39), .B(new_n685_), .C1(new_n679_), .C2(new_n686_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  NAND3_X1  g493(.A1(new_n671_), .A2(new_n274_), .A3(new_n571_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n680_), .A2(new_n682_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n274_), .B1(new_n696_), .B2(new_n571_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT41), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT41), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(new_n539_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n671_), .A2(new_n275_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n696_), .A2(new_n701_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(G22gat), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G22gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1327gat));
  INV_X1    g506(.A(new_n676_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n668_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n604_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n283_), .A3(new_n372_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n270_), .A2(new_n669_), .A3(new_n309_), .A4(new_n312_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n655_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n603_), .B2(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n536_), .A2(new_n537_), .A3(new_n519_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n537_), .B1(new_n536_), .B2(new_n519_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n565_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n489_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n572_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n601_), .A2(new_n602_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(KEYINPUT104), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n655_), .A3(new_n728_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n713_), .B(new_n714_), .C1(new_n718_), .C2(new_n729_), .ZN(new_n730_));
  AOI22_X1  g529(.A1(new_n723_), .A2(new_n724_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n731_), .B2(new_n715_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n714_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT44), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n730_), .A2(new_n734_), .A3(new_n373_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n712_), .B1(new_n735_), .B2(new_n283_), .ZN(G1328gat));
  INV_X1    g535(.A(new_n686_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n737_), .A2(G36gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n604_), .A2(new_n709_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT106), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n604_), .A2(new_n741_), .A3(new_n709_), .A4(new_n738_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n740_), .A2(new_n742_), .A3(KEYINPUT45), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT45), .B1(new_n740_), .B2(new_n742_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n730_), .A2(new_n734_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT105), .B1(new_n746_), .B2(new_n686_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n725_), .A2(new_n655_), .A3(new_n728_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n715_), .B1(new_n725_), .B2(new_n655_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n733_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n713_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n732_), .A2(KEYINPUT44), .A3(new_n733_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n751_), .A2(KEYINPUT105), .A3(new_n686_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G36gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n745_), .B1(new_n747_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT46), .B(new_n745_), .C1(new_n747_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1329gat));
  INV_X1    g558(.A(new_n571_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n288_), .B1(new_n710_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n565_), .A2(new_n288_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n746_), .B2(new_n765_), .ZN(new_n766_));
  AND4_X1   g565(.A1(new_n764_), .A2(new_n751_), .A3(new_n752_), .A4(new_n765_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT47), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n763_), .B(new_n770_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1330gat));
  NAND3_X1  g571(.A1(new_n711_), .A2(new_n286_), .A3(new_n701_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n746_), .A2(new_n701_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G50gat), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT109), .B(new_n286_), .C1(new_n746_), .C2(new_n701_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1331gat));
  NAND2_X1  g577(.A1(new_n270_), .A2(new_n312_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n677_), .A2(new_n668_), .A3(new_n308_), .A4(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G57gat), .B1(new_n780_), .B2(new_n373_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n603_), .A2(new_n309_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n779_), .A3(new_n670_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n373_), .A2(G57gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(G1332gat));
  OAI21_X1  g584(.A(G64gat), .B1(new_n780_), .B2(new_n737_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT48), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n737_), .A2(G64gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n783_), .B2(new_n788_), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n780_), .B2(new_n760_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT49), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n760_), .A2(G71gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n783_), .B2(new_n792_), .ZN(G1334gat));
  OAI21_X1  g592(.A(G78gat), .B1(new_n780_), .B2(new_n539_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n539_), .A2(G78gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT111), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n783_), .B2(new_n798_), .ZN(G1335gat));
  NAND3_X1  g598(.A1(new_n779_), .A2(new_n669_), .A3(new_n308_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n718_), .B2(new_n729_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n203_), .B1(new_n801_), .B2(new_n372_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n779_), .A2(new_n709_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n782_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(G85gat), .A3(new_n373_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT112), .Z(G1336gat));
  AOI21_X1  g606(.A(new_n204_), .B1(new_n801_), .B2(new_n686_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n804_), .A2(G92gat), .A3(new_n737_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT113), .ZN(G1337gat));
  AOI21_X1  g610(.A(new_n217_), .B1(new_n801_), .B2(new_n571_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n804_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n224_), .A2(new_n225_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n565_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n812_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n218_), .A3(new_n701_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n801_), .A2(new_n701_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G106gat), .ZN(new_n821_));
  AOI211_X1 g620(.A(KEYINPUT52), .B(new_n218_), .C1(new_n801_), .C2(new_n701_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n701_), .A2(new_n373_), .A3(new_n565_), .A4(new_n686_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n259_), .A2(new_n266_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n308_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n256_), .A2(KEYINPUT116), .A3(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n249_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(G230gat), .A3(G233gat), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n256_), .B2(KEYINPUT116), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n263_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(KEYINPUT118), .A3(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT56), .B(new_n263_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT118), .B1(new_n835_), .B2(new_n836_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n828_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n294_), .A2(new_n295_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n300_), .A2(new_n301_), .A3(new_n296_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n306_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n303_), .A2(new_n306_), .ZN(new_n845_));
  OAI22_X1  g644(.A1(new_n265_), .A2(new_n269_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n676_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n844_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n827_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n838_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n256_), .A2(KEYINPUT116), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT55), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n832_), .A3(new_n830_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n853_), .B2(new_n263_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n849_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n856_), .A2(new_n855_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n847_), .A2(KEYINPUT57), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n848_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n835_), .A2(new_n836_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n838_), .A3(new_n837_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n862_), .B1(new_n866_), .B2(new_n828_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n861_), .B1(new_n867_), .B2(new_n676_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n668_), .B1(new_n859_), .B2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT13), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT13), .B1(new_n310_), .B2(new_n311_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n308_), .A2(new_n668_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT114), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n308_), .A2(new_n875_), .A3(new_n668_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n871_), .A2(new_n872_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n870_), .B1(new_n878_), .B2(new_n717_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n874_), .A2(new_n876_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n270_), .A2(new_n880_), .A3(new_n312_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n870_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n881_), .A2(new_n655_), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n825_), .B(new_n826_), .C1(new_n869_), .C2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n847_), .B2(new_n860_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT120), .B(new_n861_), .C1(new_n867_), .C2(new_n676_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n859_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n884_), .B1(new_n889_), .B2(new_n669_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n826_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n309_), .B(new_n885_), .C1(new_n892_), .C2(new_n825_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G113gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n339_), .A3(new_n309_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1340gat));
  OAI211_X1 g695(.A(new_n779_), .B(new_n885_), .C1(new_n892_), .C2(new_n825_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G120gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n779_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n337_), .B1(new_n899_), .B2(KEYINPUT60), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n892_), .B(new_n900_), .C1(KEYINPUT60), .C2(new_n337_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n901_), .ZN(G1341gat));
  OAI211_X1 g701(.A(new_n668_), .B(new_n885_), .C1(new_n892_), .C2(new_n825_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G127gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n889_), .A2(new_n669_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n884_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n826_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n908_), .A2(G127gat), .A3(new_n669_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(new_n909_), .ZN(G1342gat));
  OAI211_X1 g709(.A(new_n655_), .B(new_n885_), .C1(new_n892_), .C2(new_n825_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G134gat), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n908_), .A2(G134gat), .A3(new_n708_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1343gat));
  NOR3_X1   g713(.A1(new_n686_), .A2(new_n571_), .A3(new_n373_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n907_), .A2(new_n701_), .A3(new_n309_), .A4(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT121), .B(G141gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1344gat));
  NOR2_X1   g717(.A1(new_n890_), .A2(new_n539_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(new_n779_), .A3(new_n915_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G148gat), .ZN(new_n921_));
  INV_X1    g720(.A(G148gat), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n919_), .A2(new_n922_), .A3(new_n779_), .A4(new_n915_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1345gat));
  NAND3_X1  g723(.A1(new_n919_), .A2(new_n668_), .A3(new_n915_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT61), .B(G155gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n926_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n919_), .A2(new_n668_), .A3(new_n915_), .A4(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1346gat));
  INV_X1    g729(.A(G162gat), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n919_), .A2(new_n931_), .A3(new_n676_), .A4(new_n915_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n919_), .A2(new_n655_), .A3(new_n915_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n931_), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n869_), .A2(new_n884_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n737_), .A2(new_n372_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n571_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n701_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n935_), .A2(new_n308_), .A3(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n941_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943_));
  INV_X1    g742(.A(G169gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n940_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n940_), .A2(new_n404_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n942_), .A2(new_n945_), .A3(new_n946_), .ZN(G1348gat));
  NOR2_X1   g746(.A1(new_n935_), .A2(new_n939_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G176gat), .B1(new_n948_), .B2(new_n779_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n701_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n899_), .A2(new_n405_), .A3(new_n937_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  NOR2_X1   g751(.A1(new_n937_), .A2(new_n669_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G183gat), .B1(new_n950_), .B2(new_n953_), .ZN(new_n954_));
  NOR4_X1   g753(.A1(new_n935_), .A2(new_n393_), .A3(new_n669_), .A4(new_n939_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT122), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n669_), .A2(new_n393_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n948_), .A2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n959_));
  INV_X1    g758(.A(new_n953_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n890_), .A2(new_n701_), .A3(new_n960_), .ZN(new_n961_));
  OAI211_X1 g760(.A(new_n958_), .B(new_n959_), .C1(G183gat), .C2(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n956_), .A2(new_n962_), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n948_), .A2(new_n676_), .A3(new_n392_), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n655_), .B(new_n938_), .C1(new_n869_), .C2(new_n884_), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n966_));
  AND3_X1   g765(.A1(new_n965_), .A2(new_n966_), .A3(G190gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n965_), .B2(G190gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n964_), .B1(new_n967_), .B2(new_n968_), .ZN(G1351gat));
  NAND2_X1  g768(.A1(new_n936_), .A2(new_n760_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n907_), .A2(new_n701_), .A3(new_n309_), .A4(new_n971_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n890_), .A2(new_n539_), .A3(new_n970_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(new_n779_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n975_), .A2(KEYINPUT124), .A3(G204gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n974_), .A2(new_n779_), .A3(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n976_), .A2(new_n978_), .ZN(G1353gat));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n980_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981_));
  AOI211_X1 g780(.A(new_n981_), .B(new_n669_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n974_), .A2(new_n982_), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n980_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n984_));
  INV_X1    g783(.A(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n983_), .A2(new_n985_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n974_), .A2(new_n984_), .A3(new_n982_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1354gat));
  NAND2_X1  g787(.A1(new_n974_), .A2(new_n676_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(KEYINPUT126), .B(G218gat), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n717_), .A2(new_n990_), .ZN(new_n991_));
  AOI22_X1  g790(.A1(new_n989_), .A2(new_n990_), .B1(new_n974_), .B2(new_n991_), .ZN(G1355gat));
endmodule


