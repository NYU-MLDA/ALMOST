//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT31), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT84), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G43gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT82), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT30), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n218_));
  OAI22_X1  g017(.A1(new_n215_), .A2(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n214_), .A2(new_n219_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G169gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n212_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n231_), .B(new_n220_), .C1(G183gat), .C2(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n232_), .A3(new_n224_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n226_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n210_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT81), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n237_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n239_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n207_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n207_), .B1(KEYINPUT84), .B2(new_n205_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G64gat), .B(G92gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(G8gat), .B(G36gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT19), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n228_), .A2(new_n232_), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n224_), .B(KEYINPUT92), .Z(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n231_), .A2(new_n220_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n216_), .A2(new_n215_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n263_), .A2(KEYINPUT91), .A3(new_n214_), .A4(new_n225_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n226_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n259_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G211gat), .A2(G218gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n270_), .B(KEYINPUT21), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G197gat), .ZN(new_n275_));
  INV_X1    g074(.A(G197gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G204gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(KEYINPUT88), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT89), .B1(new_n273_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n278_), .B2(KEYINPUT88), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n271_), .A2(new_n272_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .A4(new_n270_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n270_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n271_), .B(KEYINPUT21), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n280_), .A2(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT20), .B1(new_n267_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n234_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n256_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(new_n285_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n286_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(new_n234_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n256_), .B1(new_n267_), .B2(new_n288_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n254_), .B1(new_n292_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n299_), .A3(new_n254_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT94), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304_));
  AOI211_X1 g103(.A(KEYINPUT94), .B(new_n254_), .C1(new_n292_), .C2(new_n299_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT95), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  INV_X1    g115(.A(G141gat), .ZN(new_n317_));
  INV_X1    g116(.A(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(G155gat), .B2(G162gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n316_), .B(new_n319_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n316_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G155gat), .B(G162gat), .Z(new_n332_));
  AND3_X1   g131(.A1(new_n331_), .A2(KEYINPUT85), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT85), .B1(new_n331_), .B2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n324_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n204_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n324_), .B(new_n204_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(KEYINPUT4), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n335_), .A2(new_n340_), .A3(new_n336_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n315_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n314_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n312_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n342_), .A2(new_n312_), .A3(new_n343_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n259_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n288_), .A2(new_n226_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n290_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n256_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n289_), .A2(new_n291_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(new_n256_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n254_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT27), .A3(new_n302_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n307_), .A2(new_n347_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n335_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(KEYINPUT28), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G22gat), .B(G50gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(KEYINPUT28), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n335_), .A2(KEYINPUT29), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n296_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(G228gat), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n288_), .A2(KEYINPUT87), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n380_), .B2(new_n371_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n370_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n373_), .A2(new_n378_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n377_), .A3(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n369_), .A3(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n382_), .A2(KEYINPUT90), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT90), .B1(new_n382_), .B2(new_n385_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n368_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(KEYINPUT90), .A3(new_n385_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n249_), .A2(new_n357_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT98), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n302_), .A2(KEYINPUT94), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(new_n300_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n344_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT33), .B1(new_n344_), .B2(KEYINPUT97), .ZN(new_n398_));
  OAI22_X1  g197(.A1(new_n396_), .A2(new_n305_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n339_), .A2(new_n315_), .A3(new_n341_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n312_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n337_), .A2(new_n314_), .A3(new_n338_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n394_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n353_), .A2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n408_), .A2(new_n292_), .A3(new_n299_), .A4(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n407_), .B(new_n410_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n388_), .A2(new_n390_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n398_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n344_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n303_), .A2(new_n306_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(KEYINPUT98), .A4(new_n403_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n405_), .A2(new_n412_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n248_), .B1(new_n357_), .B2(new_n391_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n418_), .A2(KEYINPUT100), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT100), .B1(new_n418_), .B2(new_n419_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n393_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT13), .ZN(new_n423_));
  INV_X1    g222(.A(G230gat), .ZN(new_n424_));
  INV_X1    g223(.A(G233gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT10), .B(G99gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(G106gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT64), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT6), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT9), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G85gat), .A3(G92gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G85gat), .B(G92gat), .Z(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(KEYINPUT9), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n429_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT66), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT65), .B1(new_n438_), .B2(KEYINPUT7), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n431_), .B(new_n442_), .C1(new_n440_), .C2(new_n439_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT8), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT67), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(KEYINPUT67), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n443_), .A2(new_n435_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n443_), .A2(new_n435_), .A3(new_n446_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n437_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G71gat), .B(G78gat), .Z(new_n450_));
  XOR2_X1   g249(.A(G57gat), .B(G64gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT68), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G57gat), .B(G64gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT68), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n453_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n450_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n459_), .A2(new_n450_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n449_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT69), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n449_), .A2(new_n462_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT70), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n426_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n448_), .B2(new_n447_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n443_), .A2(new_n435_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n446_), .A2(new_n445_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n443_), .A2(new_n435_), .A3(new_n446_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT71), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n469_), .A2(new_n474_), .A3(new_n437_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n459_), .A2(new_n450_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n452_), .A2(new_n456_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n457_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n479_), .B2(new_n450_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n472_), .A2(new_n473_), .B1(new_n429_), .B2(new_n436_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n475_), .A2(new_n482_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n481_), .B1(new_n483_), .B2(new_n480_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n426_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n465_), .A2(KEYINPUT72), .A3(new_n481_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT5), .B(G176gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G204gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G120gat), .B(G148gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n467_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n467_), .B2(new_n490_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n423_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT13), .A3(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT75), .B(G1gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G8gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G1gat), .B(G8gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n513_), .B(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G229gat), .A3(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n512_), .A3(new_n511_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT79), .Z(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT80), .B(G113gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n518_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n502_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n422_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n475_), .A2(new_n519_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT34), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(new_n541_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n483_), .B2(new_n516_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n537_), .A2(KEYINPUT74), .A3(new_n542_), .A4(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n483_), .A2(new_n516_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n537_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT73), .B1(new_n475_), .B2(new_n519_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n543_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n549_), .A2(new_n554_), .A3(KEYINPUT36), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT37), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n567_), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT76), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n513_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n462_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT78), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n574_), .A2(new_n575_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(KEYINPUT17), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n574_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n570_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n536_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT101), .Z(new_n588_));
  INV_X1    g387(.A(new_n347_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n504_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT38), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n418_), .A2(new_n419_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT100), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n392_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n563_), .A2(new_n597_), .A3(new_n564_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n585_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n535_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n603_), .B2(new_n347_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n591_), .A2(new_n604_), .ZN(G1324gat));
  NAND2_X1  g404(.A1(new_n307_), .A2(new_n356_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n588_), .A2(new_n505_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G8gat), .B1(new_n603_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT39), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1325gat));
  OAI21_X1  g412(.A(G15gat), .B1(new_n603_), .B2(new_n249_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT41), .Z(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n588_), .A2(new_n616_), .A3(new_n248_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(new_n391_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G22gat), .B1(new_n603_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT103), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT42), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n619_), .A2(G22gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT104), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n588_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(G1327gat));
  NAND2_X1  g425(.A1(new_n565_), .A2(KEYINPUT102), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n563_), .A2(new_n597_), .A3(new_n564_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n602_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n536_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n589_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n535_), .A2(new_n585_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT105), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n422_), .A2(new_n570_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT43), .B1(new_n636_), .B2(KEYINPUT106), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n638_), .B(new_n639_), .C1(new_n422_), .C2(new_n570_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(G29gat), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT44), .B(new_n635_), .C1(new_n637_), .C2(new_n640_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n347_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n633_), .B1(new_n644_), .B2(new_n647_), .ZN(G1328gat));
  NOR3_X1   g447(.A1(new_n631_), .A2(G36gat), .A3(new_n608_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT45), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n645_), .A3(new_n606_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G36gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1329gat));
  INV_X1    g454(.A(G43gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n249_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n643_), .A2(new_n645_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n631_), .B2(new_n249_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n635_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT106), .B1(new_n596_), .B2(new_n569_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n639_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n636_), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n657_), .B1(new_n670_), .B2(KEYINPUT44), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n660_), .B1(new_n671_), .B2(new_n646_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT108), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n663_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n665_), .A2(new_n675_), .ZN(G1330gat));
  INV_X1    g475(.A(G50gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n632_), .A2(new_n677_), .A3(new_n391_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n643_), .A2(new_n645_), .A3(new_n391_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n677_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(KEYINPUT109), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n679_), .A2(new_n682_), .A3(new_n677_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n681_), .B2(new_n683_), .ZN(G1331gat));
  INV_X1    g483(.A(new_n502_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n533_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n422_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(new_n586_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n589_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n585_), .A2(new_n533_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n601_), .A2(new_n502_), .A3(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n347_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(G57gat), .B2(new_n692_), .ZN(G1332gat));
  OAI21_X1  g492(.A(G64gat), .B1(new_n691_), .B2(new_n608_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT48), .ZN(new_n695_));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n696_), .A3(new_n606_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n691_), .B2(new_n249_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT49), .ZN(new_n700_));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n688_), .A2(new_n701_), .A3(new_n248_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1334gat));
  OAI21_X1  g502(.A(G78gat), .B1(new_n691_), .B2(new_n619_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n688_), .A2(new_n707_), .A3(new_n391_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT111), .Z(G1335gat));
  AND2_X1   g509(.A1(new_n687_), .A2(new_n630_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n589_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT112), .Z(new_n713_));
  OAI211_X1 g512(.A(new_n585_), .B(new_n686_), .C1(new_n637_), .C2(new_n640_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n589_), .A2(G85gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(G1336gat));
  AOI21_X1  g516(.A(G92gat), .B1(new_n711_), .B2(new_n606_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n714_), .A2(new_n608_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g519(.A(G99gat), .B1(new_n714_), .B2(new_n249_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n249_), .A2(new_n427_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n711_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT114), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n724_), .B2(KEYINPUT51), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n726_), .B2(new_n729_), .ZN(G1338gat));
  INV_X1    g529(.A(G106gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n711_), .A2(new_n731_), .A3(new_n391_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n714_), .A2(new_n619_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G106gat), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n733_), .B(G106gat), .C1(new_n714_), .C2(new_n619_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT53), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(new_n732_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1339gat));
  NOR2_X1   g541(.A1(new_n249_), .A2(new_n391_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n606_), .A2(new_n347_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n517_), .A2(new_n523_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n520_), .A2(new_n521_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n530_), .C1(new_n747_), .C2(new_n523_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n532_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n490_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT72), .B1(new_n465_), .B2(new_n481_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n486_), .B(KEYINPUT12), .C1(new_n449_), .C2(new_n462_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n426_), .A2(KEYINPUT116), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n755_), .A2(KEYINPUT55), .A3(new_n484_), .A4(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n484_), .A2(new_n487_), .A3(KEYINPUT55), .A4(new_n489_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n756_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n752_), .A2(new_n757_), .A3(new_n760_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n494_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n494_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n496_), .B(new_n750_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n569_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT118), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n764_), .A2(new_n765_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT58), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n570_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n749_), .B1(new_n500_), .B2(new_n496_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n761_), .A2(new_n494_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n494_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n497_), .A2(new_n534_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n777_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n600_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n777_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT57), .B1(new_n629_), .B2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n770_), .A2(new_n776_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n585_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n499_), .A2(new_n501_), .A3(new_n690_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT115), .A4(new_n690_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n569_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT54), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n801_), .A3(new_n569_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n745_), .B1(new_n793_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G113gat), .B1(new_n804_), .B2(new_n533_), .ZN(new_n805_));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n533_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n785_), .B1(new_n600_), .B2(new_n784_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n629_), .A2(KEYINPUT57), .A3(new_n789_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n585_), .B1(new_n811_), .B2(new_n769_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n803_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n743_), .A4(new_n744_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n804_), .B2(new_n814_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n815_), .B(KEYINPUT119), .C1(new_n804_), .C2(new_n814_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n808_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n807_), .A2(new_n806_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n805_), .B1(new_n820_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n685_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n804_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT121), .ZN(new_n826_));
  OAI21_X1  g625(.A(G120gat), .B1(new_n816_), .B2(new_n685_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n804_), .B2(new_n602_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n818_), .A2(new_n819_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n602_), .A2(G127gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT122), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n830_), .B2(new_n832_), .ZN(G1342gat));
  AOI21_X1  g632(.A(G134gat), .B1(new_n804_), .B2(new_n600_), .ZN(new_n834_));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n570_), .ZN(G1343gat));
  INV_X1    g636(.A(new_n802_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n801_), .B1(new_n798_), .B2(new_n569_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n792_), .B2(new_n585_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n841_), .A2(new_n619_), .A3(new_n248_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n533_), .A3(new_n744_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT123), .B(G141gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1344gat));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n502_), .A3(new_n744_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n602_), .A3(new_n744_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  AND3_X1   g649(.A1(new_n842_), .A2(G162gat), .A3(new_n744_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n842_), .A2(new_n600_), .A3(new_n744_), .ZN(new_n852_));
  INV_X1    g651(.A(G162gat), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n851_), .A2(new_n570_), .B1(new_n852_), .B2(new_n853_), .ZN(G1347gat));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n608_), .A2(new_n589_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n619_), .A3(new_n248_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n812_), .B2(new_n803_), .ZN(new_n858_));
  AOI211_X1 g657(.A(KEYINPUT124), .B(new_n211_), .C1(new_n858_), .C2(new_n533_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n860_));
  INV_X1    g659(.A(new_n857_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n602_), .B1(new_n791_), .B2(new_n774_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n533_), .B(new_n861_), .C1(new_n862_), .C2(new_n840_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n863_), .B2(G169gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n855_), .B1(new_n859_), .B2(new_n864_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n534_), .B(new_n857_), .C1(new_n812_), .C2(new_n803_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n227_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT124), .B1(new_n866_), .B2(new_n211_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n860_), .A3(G169gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(KEYINPUT62), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n867_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT125), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n865_), .A2(new_n870_), .A3(new_n873_), .A4(new_n867_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1348gat));
  AOI21_X1  g674(.A(G176gat), .B1(new_n858_), .B2(new_n502_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n841_), .A2(new_n685_), .A3(new_n857_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(G176gat), .ZN(G1349gat));
  INV_X1    g677(.A(new_n858_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n879_), .A2(new_n585_), .A3(new_n261_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n841_), .A2(new_n585_), .A3(new_n857_), .ZN(new_n881_));
  INV_X1    g680(.A(G183gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n879_), .B2(new_n569_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT126), .Z(new_n885_));
  NAND3_X1  g684(.A1(new_n858_), .A2(new_n262_), .A3(new_n600_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1351gat));
  NAND3_X1  g686(.A1(new_n842_), .A2(new_n533_), .A3(new_n856_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g688(.A1(new_n842_), .A2(new_n502_), .A3(new_n856_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT127), .B(G204gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1353gat));
  NAND3_X1  g691(.A1(new_n842_), .A2(new_n602_), .A3(new_n856_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n893_), .B2(new_n895_), .ZN(G1354gat));
  AND3_X1   g695(.A1(new_n842_), .A2(G218gat), .A3(new_n856_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n842_), .A2(new_n600_), .A3(new_n856_), .ZN(new_n898_));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n570_), .B1(new_n898_), .B2(new_n899_), .ZN(G1355gat));
endmodule


