//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G169gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .A4(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT82), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n214_), .B(new_n213_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(new_n212_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n211_), .B(new_n217_), .C1(KEYINPUT82), .C2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n218_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G183gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n224_), .B2(G183gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n223_), .A2(new_n225_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n233_), .B2(new_n210_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n222_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n221_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n236_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT31), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT31), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n245_), .A2(KEYINPUT83), .A3(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n241_), .B(new_n247_), .Z(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G43gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n248_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G22gat), .B(G50gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n257_));
  AND2_X1   g056(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G141gat), .ZN(new_n260_));
  INV_X1    g059(.A(G148gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT85), .ZN(new_n262_));
  INV_X1    g061(.A(new_n254_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n262_), .A2(KEYINPUT3), .B1(new_n263_), .B2(KEYINPUT2), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n259_), .B(new_n264_), .C1(KEYINPUT3), .C2(new_n262_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G155gat), .B(G162gat), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n261_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n269_), .A2(new_n256_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT87), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT87), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n267_), .A2(new_n275_), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n253_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(new_n280_), .A3(new_n252_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n279_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT88), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(KEYINPUT88), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n289_), .A2(new_n290_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n291_), .B(KEYINPUT21), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n296_), .A2(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(G228gat), .B(G233gat), .C1(new_n287_), .C2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n277_), .A2(new_n279_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n297_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n301_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G78gat), .B(G106gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT90), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n312_));
  INV_X1    g111(.A(new_n309_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n286_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n316_), .A3(new_n309_), .ZN(new_n317_));
  OAI221_X1 g116(.A(new_n301_), .B1(KEYINPUT91), .B2(new_n313_), .C1(new_n302_), .C2(new_n307_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n285_), .A3(new_n283_), .A4(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT97), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n274_), .A2(new_n321_), .A3(new_n276_), .A4(new_n244_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n274_), .A2(new_n276_), .A3(new_n244_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT97), .B1(new_n273_), .B2(new_n244_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT4), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n274_), .A2(new_n327_), .A3(new_n276_), .A4(new_n244_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT99), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT98), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n331_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G85gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT0), .B(G57gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT33), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT20), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n305_), .B2(new_n236_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n218_), .B1(new_n223_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n234_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n203_), .A2(new_n208_), .A3(new_n205_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n210_), .B(KEYINPUT93), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n219_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT94), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n300_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n347_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n347_), .A2(KEYINPUT95), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G8gat), .B(G36gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n356_), .A2(new_n350_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n305_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n300_), .A2(new_n221_), .A3(new_n235_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT20), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n344_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n362_), .A2(new_n368_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n360_), .A2(new_n361_), .B1(new_n344_), .B2(new_n372_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n368_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n333_), .A2(KEYINPUT33), .A3(new_n334_), .A4(new_n338_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n326_), .A2(new_n331_), .A3(new_n330_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n338_), .B1(new_n325_), .B2(new_n332_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n341_), .A2(new_n378_), .A3(new_n379_), .A4(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n370_), .A2(KEYINPUT20), .A3(new_n345_), .A4(new_n371_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n305_), .B2(new_n236_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n300_), .B(new_n350_), .C1(new_n219_), .C2(new_n353_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n345_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n391_), .B2(new_n376_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n339_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n338_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n320_), .B1(new_n383_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n395_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n320_), .A2(new_n398_), .A3(new_n339_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n374_), .A2(KEYINPUT102), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n367_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(KEYINPUT101), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT101), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n367_), .C1(new_n385_), .C2(new_n389_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT102), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n376_), .A2(new_n406_), .A3(new_n368_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n400_), .A2(new_n403_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n401_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n399_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n251_), .B1(new_n397_), .B2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n410_), .A2(new_n320_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n398_), .A2(new_n339_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(new_n251_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G29gat), .B(G36gat), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n418_), .A2(KEYINPUT74), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(KEYINPUT74), .ZN(new_n420_));
  XOR2_X1   g219(.A(G43gat), .B(G50gat), .Z(new_n421_));
  OR3_X1    g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT15), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G22gat), .ZN(new_n427_));
  INV_X1    g226(.A(G1gat), .ZN(new_n428_));
  INV_X1    g227(.A(G8gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G1gat), .B(G8gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT15), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n426_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n433_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G229gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n422_), .A2(new_n433_), .A3(new_n423_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(new_n441_), .B2(new_n436_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G113gat), .B(G141gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G169gat), .B(G197gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n447_), .B(new_n445_), .C1(new_n440_), .C2(new_n442_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n452_), .B(KEYINPUT79), .Z(new_n453_));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G232gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT34), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT35), .Z(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(KEYINPUT6), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT10), .B(G99gat), .Z(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(KEYINPUT65), .A3(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT67), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n474_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n475_));
  AND3_X1   g274(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n472_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n473_), .B1(new_n472_), .B2(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n465_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI22_X1  g280(.A1(KEYINPUT68), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n482_), .B(new_n485_), .C1(new_n459_), .C2(new_n461_), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n489_), .A2(new_n466_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT69), .A3(new_n466_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n486_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n426_), .A2(new_n434_), .B1(new_n481_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n481_), .A2(new_n496_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n424_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT75), .B(new_n457_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n497_), .A2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n456_), .A2(KEYINPUT35), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT75), .B1(new_n501_), .B2(new_n457_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n454_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G190gat), .B(G218gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(G134gat), .B(G162gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n509_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n505_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  OAI221_X1 g313(.A(new_n454_), .B1(new_n514_), .B2(new_n510_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(KEYINPUT37), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT37), .B1(new_n513_), .B2(new_n515_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT71), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n464_), .A2(new_n463_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT65), .B1(new_n466_), .B2(new_n467_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n471_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n478_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT67), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n472_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n523_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n485_), .A2(new_n482_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n490_), .B1(new_n462_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n493_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n486_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n521_), .B1(new_n529_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n481_), .A2(new_n496_), .A3(new_n520_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G57gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(G64gat), .ZN(new_n542_));
  INV_X1    g341(.A(G64gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(G57gat), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT70), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT11), .B1(new_n540_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G71gat), .B(G78gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(new_n539_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT70), .B1(new_n542_), .B2(new_n544_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT11), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT11), .B(new_n547_), .C1(new_n540_), .C2(new_n545_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n536_), .A2(new_n537_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n498_), .A2(new_n558_), .A3(KEYINPUT12), .A4(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT64), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT72), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n565_));
  AOI211_X1 g364(.A(new_n565_), .B(new_n562_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n498_), .B2(new_n555_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n498_), .B2(new_n555_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G120gat), .B(G148gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n569_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G127gat), .B(G155gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT17), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n585_), .A2(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n433_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n556_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n592_));
  AOI211_X1 g391(.A(new_n587_), .B(new_n588_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n591_), .A2(KEYINPUT71), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(KEYINPUT71), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n587_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n576_), .A2(KEYINPUT13), .A3(new_n578_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n581_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n519_), .A2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n417_), .A2(new_n453_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n428_), .A3(new_n414_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n513_), .A2(new_n515_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n581_), .A2(new_n599_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n452_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n598_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n414_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n605_), .A2(new_n606_), .A3(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n602_), .A2(new_n429_), .A3(new_n410_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  INV_X1    g417(.A(new_n613_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n410_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n620_), .B2(G8gat), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT39), .B(new_n429_), .C1(new_n619_), .C2(new_n410_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n617_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n613_), .B2(new_n251_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  INV_X1    g425(.A(new_n251_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n602_), .A2(new_n238_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(new_n320_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G22gat), .B1(new_n613_), .B2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n602_), .A2(new_n634_), .A3(new_n320_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1327gat));
  NOR3_X1   g435(.A1(new_n609_), .A2(new_n610_), .A3(new_n598_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n417_), .B2(new_n519_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n518_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n516_), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT43), .B(new_n641_), .C1(new_n412_), .C2(new_n416_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n637_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT44), .B(new_n637_), .C1(new_n639_), .C2(new_n642_), .ZN(new_n646_));
  AND4_X1   g445(.A1(G29gat), .A2(new_n645_), .A3(new_n414_), .A4(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n607_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n609_), .A2(new_n648_), .A3(new_n598_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n417_), .A2(new_n453_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n414_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n647_), .A2(new_n652_), .ZN(G1328gat));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n656_));
  INV_X1    g455(.A(G36gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n410_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n656_), .B1(new_n651_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n656_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n650_), .A2(new_n661_), .A3(new_n658_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n645_), .A2(new_n410_), .A3(new_n646_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(G36gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1329gat));
  NAND4_X1  g466(.A1(new_n645_), .A2(G43gat), .A3(new_n627_), .A4(new_n646_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n650_), .A2(new_n251_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(G43gat), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g470(.A1(G50gat), .A2(new_n645_), .A3(new_n320_), .A4(new_n646_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G50gat), .B1(new_n651_), .B2(new_n320_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1331gat));
  INV_X1    g473(.A(new_n453_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n609_), .A2(new_n598_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n608_), .A2(new_n675_), .A3(new_n677_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT107), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT107), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n614_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n452_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(new_n641_), .A3(new_n677_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n541_), .A3(new_n414_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1332gat));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n543_), .A3(new_n410_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT48), .ZN(new_n688_));
  INV_X1    g487(.A(new_n681_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n410_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(G64gat), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT48), .B(new_n543_), .C1(new_n689_), .C2(new_n410_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n684_), .A2(new_n694_), .A3(new_n627_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G71gat), .B1(new_n681_), .B2(new_n251_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(G1334gat));
  NOR2_X1   g498(.A1(new_n630_), .A2(G78gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT108), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n684_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G78gat), .B1(new_n681_), .B2(new_n630_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT50), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT50), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(G1335gat));
  INV_X1    g505(.A(new_n609_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(new_n648_), .A3(new_n598_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n683_), .A2(KEYINPUT109), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT109), .B1(new_n683_), .B2(new_n708_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n487_), .A3(new_n414_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n639_), .A2(new_n642_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT110), .Z(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n414_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n713_), .B1(new_n720_), .B2(new_n487_), .ZN(G1336gat));
  NAND3_X1  g520(.A1(new_n712_), .A2(new_n488_), .A3(new_n410_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n410_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n488_), .ZN(G1337gat));
  OAI21_X1  g524(.A(G99gat), .B1(new_n717_), .B2(new_n251_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n627_), .A2(new_n464_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n711_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT51), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n726_), .B(new_n730_), .C1(new_n711_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1338gat));
  OAI211_X1 g531(.A(new_n320_), .B(new_n716_), .C1(new_n639_), .C2(new_n642_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(G106gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n733_), .B2(G106gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n738_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n712_), .A2(new_n463_), .A3(new_n320_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT53), .B1(new_n739_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n737_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT52), .A3(new_n735_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(G1339gat));
  INV_X1    g547(.A(KEYINPUT57), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n607_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n436_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n435_), .A2(new_n751_), .A3(new_n438_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n445_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n441_), .A2(new_n436_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n752_), .B(new_n753_), .C1(new_n754_), .C2(new_n438_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n446_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n579_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n452_), .A2(new_n578_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n557_), .A2(new_n562_), .A3(new_n559_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n560_), .A2(new_n563_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n567_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(new_n577_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n565_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n562_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT72), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n769_), .A3(new_n764_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n760_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(KEYINPUT55), .B2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n758_), .B1(new_n766_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n757_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT113), .B(new_n758_), .C1(new_n766_), .C2(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n750_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT115), .ZN(new_n780_));
  INV_X1    g579(.A(new_n758_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n575_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n759_), .B(new_n577_), .C1(new_n770_), .C2(new_n772_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT113), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n766_), .A2(new_n774_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n776_), .A3(new_n781_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(new_n757_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n750_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT114), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n578_), .B(new_n756_), .C1(new_n766_), .C2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n578_), .A2(new_n756_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n782_), .B2(KEYINPUT114), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(KEYINPUT58), .C1(KEYINPUT114), .C2(new_n786_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n519_), .A3(new_n799_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n784_), .A2(KEYINPUT113), .B1(new_n579_), .B2(new_n756_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n607_), .B1(new_n801_), .B2(new_n787_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(KEYINPUT57), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n611_), .B1(new_n791_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n601_), .B2(new_n675_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n519_), .A2(new_n600_), .A3(KEYINPUT54), .A4(new_n453_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n804_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n413_), .A2(new_n414_), .A3(new_n627_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(KEYINPUT59), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n648_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n749_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(new_n780_), .A3(new_n800_), .A4(new_n790_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n808_), .B1(new_n817_), .B2(new_n611_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n818_), .B2(new_n811_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n813_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820_), .B2(new_n675_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n810_), .A2(KEYINPUT116), .A3(new_n812_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n818_), .B2(new_n811_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n452_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n827_), .ZN(G1340gat));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n829_), .A2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n822_), .A2(new_n824_), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n707_), .B1(new_n813_), .B2(new_n819_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n829_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT117), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n832_), .B(new_n836_), .C1(new_n833_), .C2(new_n829_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n820_), .B2(new_n611_), .ZN(new_n839_));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n825_), .A2(new_n840_), .A3(new_n598_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1342gat));
  OAI21_X1  g641(.A(G134gat), .B1(new_n820_), .B2(new_n641_), .ZN(new_n843_));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n825_), .A2(new_n844_), .A3(new_n607_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1343gat));
  NAND3_X1  g645(.A1(new_n414_), .A2(new_n320_), .A3(new_n251_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n818_), .A2(new_n410_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n452_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n609_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n598_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(G162gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n848_), .A2(new_n856_), .A3(new_n607_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n848_), .A2(new_n519_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1347gat));
  NAND2_X1  g658(.A1(new_n415_), .A2(new_n410_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT118), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n861_), .A2(new_n630_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n810_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n610_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n207_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n203_), .A3(new_n208_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(G1348gat));
  INV_X1    g668(.A(new_n863_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G176gat), .B1(new_n870_), .B2(new_n609_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n810_), .A2(KEYINPUT119), .A3(new_n630_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n818_), .B2(new_n320_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n872_), .A2(new_n874_), .A3(new_n861_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n707_), .A2(new_n205_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n871_), .B1(new_n875_), .B2(new_n876_), .ZN(G1349gat));
  NOR3_X1   g676(.A1(new_n863_), .A2(new_n348_), .A3(new_n611_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n598_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n226_), .ZN(G1350gat));
  NAND2_X1  g679(.A1(new_n607_), .A2(new_n223_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT121), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n870_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n810_), .A2(new_n519_), .A3(new_n862_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n884_), .A2(KEYINPUT120), .A3(G190gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT120), .B1(new_n884_), .B2(G190gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT122), .B(new_n883_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1351gat));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  INV_X1    g691(.A(new_n399_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n410_), .A3(new_n251_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n892_), .B1(new_n810_), .B2(new_n895_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n818_), .A2(KEYINPUT123), .A3(new_n894_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n452_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(G197gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(KEYINPUT125), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT123), .B1(new_n818_), .B2(new_n894_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n750_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT115), .B(new_n903_), .C1(new_n801_), .C2(new_n787_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n789_), .B1(new_n788_), .B2(new_n750_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n798_), .B1(new_n786_), .B2(KEYINPUT114), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n641_), .B1(new_n907_), .B2(new_n792_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n799_), .A2(new_n908_), .B1(new_n815_), .B2(new_n749_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n598_), .B1(new_n906_), .B2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n892_), .B(new_n895_), .C1(new_n910_), .C2(new_n808_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n610_), .B1(new_n902_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n901_), .B1(new_n912_), .B2(G197gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n900_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n902_), .A2(new_n911_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n610_), .A2(new_n899_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n917_), .ZN(new_n919_));
  AOI211_X1 g718(.A(KEYINPUT124), .B(new_n919_), .C1(new_n902_), .C2(new_n911_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n914_), .A2(new_n921_), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n609_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g723(.A(new_n611_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n916_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT126), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n926_), .B(new_n928_), .ZN(G1354gat));
  AND2_X1   g728(.A1(new_n519_), .A2(G218gat), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n916_), .A2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n648_), .B1(new_n902_), .B2(new_n911_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(G218gat), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n931_), .B(KEYINPUT127), .C1(G218gat), .C2(new_n932_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1355gat));
endmodule


