//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  AND2_X1   g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT65), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT7), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n211_), .A2(new_n206_), .A3(new_n207_), .A4(KEYINPUT65), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n213_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n210_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT8), .B(new_n205_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n209_), .A2(new_n218_), .A3(new_n212_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n205_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(G92gat), .ZN(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n204_), .B1(new_n203_), .B2(KEYINPUT9), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT10), .B(G99gat), .Z(new_n234_));
  AOI22_X1  g033(.A1(new_n234_), .A2(new_n207_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n226_), .A2(new_n227_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n224_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G78gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n239_), .B(new_n240_), .C1(KEYINPUT11), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G64gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G57gat), .ZN(new_n244_));
  INV_X1    g043(.A(G57gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G64gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT11), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n247_), .B2(new_n238_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n242_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n237_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n237_), .A2(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n237_), .A2(new_n252_), .A3(KEYINPUT12), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n237_), .A2(new_n252_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n237_), .A2(new_n252_), .ZN(new_n261_));
  OAI211_X1 g060(.A(G230gat), .B(G233gat), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G120gat), .B(G148gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(G176gat), .B(G204gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT70), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n259_), .A2(new_n262_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n202_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n259_), .A2(new_n262_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n268_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n259_), .A2(new_n262_), .A3(new_n269_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT71), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT13), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT72), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n270_), .A2(new_n271_), .A3(new_n202_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT71), .B1(new_n274_), .B2(new_n275_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT13), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT73), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT105), .ZN(new_n290_));
  INV_X1    g089(.A(G155gat), .ZN(new_n291_));
  INV_X1    g090(.A(G162gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT92), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT92), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT95), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  INV_X1    g102(.A(G141gat), .ZN(new_n304_));
  INV_X1    g103(.A(G148gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  OAI22_X1  g106(.A1(KEYINPUT95), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n295_), .B1(new_n301_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT96), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT96), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n312_), .B(new_n295_), .C1(new_n301_), .C2(new_n309_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT93), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n294_), .A2(new_n315_), .A3(KEYINPUT1), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n293_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n294_), .B2(KEYINPUT1), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT94), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n294_), .A2(KEYINPUT1), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT93), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT94), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n293_), .A4(new_n316_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n294_), .A2(KEYINPUT1), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n297_), .A2(new_n299_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n314_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G120gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n311_), .A2(new_n313_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT0), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT102), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  AND3_X1   g143(.A1(new_n314_), .A2(new_n332_), .A3(new_n328_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n332_), .B1(new_n314_), .B2(new_n328_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n329_), .A2(new_n347_), .A3(new_n333_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n337_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n338_), .B(new_n344_), .C1(new_n348_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT103), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT33), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n352_), .B(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n334_), .A2(KEYINPUT4), .A3(new_n336_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n337_), .A3(new_n349_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n334_), .A2(new_n336_), .A3(new_n350_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT104), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n342_), .B(new_n343_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n357_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n368_), .A2(KEYINPUT21), .ZN(new_n369_));
  XOR2_X1   g168(.A(G197gat), .B(G204gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(KEYINPUT21), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n370_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G190gat), .ZN(new_n377_));
  INV_X1    g176(.A(G183gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT25), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G183gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n376_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(G183gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n378_), .A2(KEYINPUT25), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT86), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(KEYINPUT87), .A3(new_n377_), .A4(new_n381_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(KEYINPUT24), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT88), .A3(KEYINPUT23), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G183gat), .A3(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT88), .B1(new_n398_), .B2(KEYINPUT23), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n395_), .B(new_n397_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n391_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G169gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT22), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT22), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G169gat), .ZN(new_n410_));
  INV_X1    g209(.A(G176gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n394_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n398_), .A2(KEYINPUT23), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT89), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n398_), .A2(new_n416_), .A3(KEYINPUT23), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n417_), .A3(new_n401_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G183gat), .A2(G190gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n413_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n375_), .B1(new_n406_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT25), .B(G183gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n425_));
  NOR2_X1   g224(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n424_), .A2(new_n377_), .B1(new_n427_), .B2(new_n392_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT100), .B1(new_n429_), .B2(new_n394_), .ZN(new_n430_));
  OAI211_X1 g229(.A(KEYINPUT100), .B(new_n394_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n393_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n428_), .B(new_n418_), .C1(new_n430_), .C2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n420_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n412_), .A2(KEYINPUT101), .A3(new_n394_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT101), .B1(new_n412_), .B2(new_n394_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n372_), .A2(new_n374_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT20), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n367_), .B1(new_n423_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n406_), .B2(new_n422_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n438_), .A2(new_n375_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT20), .B(new_n366_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT18), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n441_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n363_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n290_), .B1(new_n355_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT108), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n352_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n356_), .A2(new_n350_), .A3(new_n349_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n456_), .A2(KEYINPUT108), .A3(new_n338_), .A4(new_n344_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n338_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n360_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n441_), .A2(new_n444_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n448_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n442_), .B2(new_n443_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n366_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT107), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT106), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n432_), .A2(new_n430_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n427_), .A2(new_n392_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n424_), .A2(new_n377_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n418_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT101), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n413_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n412_), .A2(KEYINPUT101), .A3(new_n394_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n403_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n401_), .A3(new_n399_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n475_), .A2(new_n476_), .B1(new_n478_), .B2(new_n420_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n468_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n433_), .A2(new_n437_), .A3(KEYINPUT106), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n439_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n467_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n423_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n433_), .A2(new_n437_), .A3(KEYINPUT106), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT106), .B1(new_n433_), .B2(new_n437_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n375_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT107), .A3(KEYINPUT20), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n466_), .B1(new_n490_), .B2(new_n366_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n460_), .B(new_n464_), .C1(new_n491_), .C2(new_n463_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n352_), .B1(new_n353_), .B2(KEYINPUT33), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n456_), .A2(new_n338_), .A3(new_n344_), .A4(new_n354_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n495_), .A2(KEYINPUT105), .A3(new_n451_), .A4(new_n363_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n453_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n335_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT28), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G228gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT97), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n498_), .B1(new_n314_), .B2(new_n328_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n375_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n439_), .B(new_n503_), .C1(new_n335_), .C2(new_n498_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G22gat), .B(G50gat), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n508_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n313_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n516_), .A2(new_n306_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n312_), .B1(new_n517_), .B2(new_n295_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n325_), .A2(new_n327_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT29), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n503_), .B1(new_n521_), .B2(new_n439_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n507_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n514_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n511_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n501_), .B1(new_n513_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n512_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n525_), .A3(new_n511_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n500_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n406_), .A2(KEYINPUT30), .A3(new_n422_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G227gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G15gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT90), .ZN(new_n534_));
  INV_X1    g333(.A(G15gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n532_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G71gat), .B(G99gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G43gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n540_), .A2(G43gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(G43gat), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n534_), .A2(new_n538_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n404_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n421_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n531_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT91), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n531_), .A2(new_n546_), .A3(new_n549_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n546_), .B1(new_n531_), .B2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT31), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n556_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n332_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n562_));
  AOI211_X1 g361(.A(KEYINPUT31), .B(new_n555_), .C1(new_n551_), .C2(new_n553_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n333_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n527_), .A2(new_n530_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n497_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n528_), .A2(new_n500_), .A3(new_n529_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n500_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n561_), .B(new_n564_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(new_n564_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n460_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n451_), .A2(KEYINPUT27), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n480_), .A2(new_n481_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n483_), .B1(new_n576_), .B2(new_n375_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n423_), .B1(new_n577_), .B2(KEYINPUT107), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n367_), .B1(new_n578_), .B2(new_n484_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n448_), .B1(new_n579_), .B2(new_n466_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT27), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n450_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT109), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT109), .B(new_n582_), .C1(new_n491_), .C2(new_n462_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n573_), .B(new_n575_), .C1(new_n583_), .C2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n566_), .B1(new_n572_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT82), .B(G8gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G1gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT14), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G1gat), .B(G8gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G29gat), .B(G36gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G43gat), .B(G50gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n595_), .B(new_n598_), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(KEYINPUT15), .ZN(new_n600_));
  MUX2_X1   g399(.A(new_n600_), .B(new_n598_), .S(new_n595_), .Z(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  MUX2_X1   g401(.A(new_n599_), .B(new_n601_), .S(new_n602_), .Z(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G169gat), .B(G197gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT85), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n603_), .B(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n224_), .A2(new_n236_), .A3(new_n598_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT75), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n224_), .A2(new_n236_), .A3(new_n611_), .A4(new_n598_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n237_), .B2(new_n600_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT76), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n620_), .A2(KEYINPUT76), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n613_), .A2(new_n622_), .A3(new_n618_), .A4(new_n621_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT77), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT36), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n627_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(KEYINPUT79), .A2(KEYINPUT80), .A3(KEYINPUT37), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT79), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n627_), .A2(new_n637_), .A3(new_n628_), .A4(new_n633_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT78), .Z(new_n642_));
  AOI211_X1 g441(.A(new_n623_), .B(new_n625_), .C1(new_n613_), .C2(new_n618_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n628_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT81), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(KEYINPUT80), .A3(new_n634_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(new_n646_), .B2(new_n650_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n595_), .B(new_n252_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(G231gat), .A2(G233gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT83), .Z(new_n656_));
  XNOR2_X1  g455(.A(new_n654_), .B(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(G127gat), .B(G155gat), .Z(new_n658_));
  XNOR2_X1  g457(.A(G183gat), .B(G211gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT17), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n657_), .A2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n662_), .A2(KEYINPUT17), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n653_), .A2(new_n668_), .ZN(new_n669_));
  AND4_X1   g468(.A1(new_n289_), .A2(new_n587_), .A3(new_n608_), .A4(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n590_), .A3(new_n460_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT112), .Z(new_n674_));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n489_), .A2(new_n485_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT107), .B1(new_n488_), .B2(KEYINPUT20), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n366_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n466_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n462_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n582_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n675_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n460_), .B(new_n574_), .C1(new_n682_), .C2(new_n584_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n569_), .A2(new_n571_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n683_), .A2(new_n684_), .B1(new_n497_), .B2(new_n565_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n645_), .A2(new_n634_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT111), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n280_), .A2(new_n286_), .A3(new_n608_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n280_), .A2(new_n286_), .A3(KEYINPUT110), .A4(new_n608_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n668_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G1gat), .B1(new_n695_), .B2(new_n573_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n674_), .B(new_n696_), .C1(new_n672_), .C2(new_n671_), .ZN(G1324gat));
  NAND2_X1  g496(.A1(new_n682_), .A2(new_n584_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n575_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n670_), .A2(new_n699_), .A3(new_n589_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n689_), .A2(new_n699_), .A3(new_n694_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT39), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G8gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G8gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g505(.A(G15gat), .B1(new_n695_), .B2(new_n570_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n708_));
  OR2_X1    g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n570_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n670_), .A2(new_n535_), .A3(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n710_), .A3(new_n712_), .ZN(G1326gat));
  INV_X1    g512(.A(G22gat), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n567_), .A2(new_n568_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n670_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n717_));
  INV_X1    g516(.A(new_n695_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n715_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(G22gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT42), .B(new_n714_), .C1(new_n718_), .C2(new_n715_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n720_), .B2(new_n721_), .ZN(G1327gat));
  NAND2_X1  g521(.A1(new_n668_), .A2(new_n687_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n685_), .A2(new_n690_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(new_n460_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n667_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n648_), .A2(new_n649_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n627_), .A2(new_n628_), .ZN(new_n728_));
  AOI22_X1  g527(.A1(new_n636_), .A2(new_n638_), .B1(new_n728_), .B2(new_n642_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT81), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n685_), .A2(KEYINPUT43), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n587_), .B2(new_n653_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n726_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n738_), .A2(G29gat), .A3(new_n460_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n726_), .B(KEYINPUT44), .C1(new_n733_), .C2(new_n735_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n725_), .B1(new_n739_), .B2(new_n740_), .ZN(G1328gat));
  NAND2_X1  g540(.A1(KEYINPUT116), .A2(KEYINPUT46), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n699_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G36gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT114), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n747_), .A3(G36gat), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(KEYINPUT116), .A2(KEYINPUT46), .ZN(new_n750_));
  INV_X1    g549(.A(G36gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n724_), .A2(new_n751_), .A3(new_n699_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n753_));
  OR2_X1    g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n753_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n743_), .B1(new_n749_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n699_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT114), .B(new_n751_), .C1(new_n759_), .C2(new_n740_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n747_), .B1(new_n744_), .B2(G36gat), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n743_), .B(new_n756_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n742_), .B1(new_n757_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n756_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT117), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(KEYINPUT116), .A3(KEYINPUT46), .A4(new_n762_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(G1329gat));
  NAND4_X1  g567(.A1(new_n738_), .A2(G43gat), .A3(new_n711_), .A4(new_n740_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n724_), .A2(new_n711_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(G43gat), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g571(.A(G50gat), .B1(new_n724_), .B2(new_n715_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n738_), .A2(G50gat), .A3(new_n715_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n740_), .ZN(G1331gat));
  INV_X1    g574(.A(new_n287_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n608_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n777_), .A2(new_n669_), .A3(new_n587_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n245_), .A3(new_n460_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n608_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n667_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n289_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n689_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n460_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n779_), .B1(new_n784_), .B2(new_n245_), .ZN(G1332gat));
  NAND3_X1  g584(.A1(new_n778_), .A2(new_n243_), .A3(new_n699_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n699_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G64gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT48), .B(new_n243_), .C1(new_n783_), .C2(new_n699_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT118), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n783_), .B2(new_n711_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT49), .Z(new_n795_));
  NAND3_X1  g594(.A1(new_n778_), .A2(new_n793_), .A3(new_n711_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1334gat));
  INV_X1    g596(.A(G78gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n783_), .B2(new_n715_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT50), .Z(new_n800_));
  NAND3_X1  g599(.A1(new_n778_), .A2(new_n798_), .A3(new_n715_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1335gat));
  OR2_X1    g601(.A1(new_n733_), .A2(new_n735_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n668_), .A3(new_n777_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n573_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n685_), .A2(new_n608_), .A3(new_n723_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n288_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n230_), .A3(new_n460_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n805_), .A2(new_n809_), .ZN(G1336gat));
  AOI21_X1  g609(.A(G92gat), .B1(new_n808_), .B2(new_n699_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n803_), .A2(new_n668_), .A3(new_n777_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n758_), .A2(new_n229_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n804_), .B2(new_n570_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n711_), .A2(new_n234_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n807_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g617(.A(new_n207_), .B1(new_n812_), .B2(new_n715_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(KEYINPUT119), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  INV_X1    g621(.A(new_n715_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G106gat), .B1(new_n804_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n824_), .B2(KEYINPUT52), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT52), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n821_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n808_), .A2(new_n207_), .A3(new_n715_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT53), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1339gat));
  AND3_X1   g632(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT55), .A3(new_n257_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n259_), .A2(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n837_), .C1(new_n257_), .C2(new_n834_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n838_), .A2(KEYINPUT56), .A3(new_n268_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n838_), .B2(new_n268_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n275_), .B(new_n608_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n599_), .B1(G229gat), .B2(G233gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n601_), .A2(new_n602_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n606_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n846_), .A2(new_n276_), .A3(new_n272_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n686_), .B1(new_n842_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n849_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n839_), .A2(new_n840_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n270_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT58), .B1(new_n853_), .B2(new_n846_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n846_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n653_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n850_), .B(new_n851_), .C1(new_n854_), .C2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n668_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n781_), .A2(new_n279_), .A3(new_n278_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n732_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT54), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n699_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT59), .ZN(new_n865_));
  OAI21_X1  g664(.A(G113gat), .B1(new_n865_), .B2(new_n780_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n780_), .A2(G113gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n864_), .B2(new_n867_), .ZN(G1340gat));
  OAI21_X1  g667(.A(G120gat), .B1(new_n865_), .B2(new_n289_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n864_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n287_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n869_), .A2(new_n875_), .ZN(G1341gat));
  OAI21_X1  g675(.A(G127gat), .B1(new_n865_), .B2(new_n668_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n668_), .A2(G127gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n864_), .B2(new_n878_), .ZN(G1342gat));
  OAI21_X1  g678(.A(G134gat), .B1(new_n865_), .B2(new_n732_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n864_), .A2(G134gat), .A3(new_n686_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1343gat));
  INV_X1    g681(.A(new_n861_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n668_), .B2(new_n857_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n571_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n460_), .A3(new_n758_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n780_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n304_), .ZN(G1344gat));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n289_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n305_), .ZN(G1345gat));
  NOR2_X1   g689(.A1(new_n886_), .A2(new_n668_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT61), .B(G155gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n886_), .B2(new_n732_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n687_), .A2(new_n292_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n886_), .B2(new_n895_), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n408_), .A2(new_n410_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n758_), .A2(new_n570_), .A3(new_n460_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n608_), .ZN(new_n899_));
  OR4_X1    g698(.A1(new_n897_), .A2(new_n884_), .A3(new_n715_), .A4(new_n899_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n899_), .B(KEYINPUT121), .Z(new_n901_));
  NAND3_X1  g700(.A1(new_n862_), .A2(new_n823_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n862_), .A2(KEYINPUT122), .A3(new_n901_), .A4(new_n823_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(G169gat), .A3(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n900_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n862_), .A2(new_n823_), .A3(new_n898_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n411_), .B1(new_n910_), .B2(new_n776_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n912_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT124), .B1(new_n884_), .B2(new_n715_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n862_), .A2(new_n916_), .A3(new_n823_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n898_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n289_), .A2(new_n411_), .A3(new_n919_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n913_), .A2(new_n914_), .B1(new_n918_), .B2(new_n920_), .ZN(G1349gat));
  NOR3_X1   g720(.A1(new_n910_), .A2(new_n424_), .A3(new_n668_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n919_), .A2(new_n668_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n915_), .A2(new_n917_), .A3(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(KEYINPUT125), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(G183gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(KEYINPUT125), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n922_), .B1(new_n926_), .B2(new_n927_), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n910_), .B2(new_n732_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n687_), .A2(new_n377_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n910_), .B2(new_n930_), .ZN(G1351gat));
  NOR2_X1   g730(.A1(new_n758_), .A2(new_n460_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n885_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n780_), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT126), .B(G197gat), .Z(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1352gat));
  INV_X1    g735(.A(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n288_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g738(.A1(new_n933_), .A2(new_n668_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AND2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n940_), .B2(new_n941_), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n937_), .B2(new_n687_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n653_), .A2(G218gat), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n946_), .B(KEYINPUT127), .Z(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n937_), .B2(new_n947_), .ZN(G1355gat));
endmodule


