//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT86), .B1(new_n207_), .B2(KEYINPUT85), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(new_n209_), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n208_), .A2(new_n209_), .B1(new_n212_), .B2(new_n207_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n206_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n207_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(new_n204_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT1), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n218_), .B(new_n219_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(new_n227_), .A3(new_n223_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(KEYINPUT4), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT95), .B(KEYINPUT4), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n230_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n233_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n231_), .A2(new_n235_), .B1(new_n237_), .B2(new_n232_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n231_), .A2(new_n235_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n237_), .A2(new_n232_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT99), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT99), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n238_), .A2(new_n250_), .A3(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT19), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  INV_X1    g055(.A(G197gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT88), .B1(new_n257_), .B2(G204gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G197gat), .B(G204gat), .Z(new_n262_));
  NAND4_X1  g061(.A1(new_n262_), .A2(KEYINPUT21), .A3(new_n256_), .A4(new_n258_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n256_), .A2(KEYINPUT21), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT22), .B(G169gat), .Z(new_n269_));
  INV_X1    g068(.A(KEYINPUT81), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT23), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  OAI221_X1 g078(.A(new_n268_), .B1(G176gat), .B2(new_n269_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT25), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G183gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(KEYINPUT24), .A3(new_n268_), .A4(new_n291_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n272_), .A2(new_n276_), .A3(new_n274_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n276_), .A2(new_n271_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n294_), .B(new_n299_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n280_), .B1(new_n289_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n267_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT26), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(KEYINPUT78), .A3(G190gat), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n306_), .A2(new_n308_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n294_), .A2(new_n309_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n299_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n290_), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n313_), .A2(new_n298_), .A3(KEYINPUT80), .A4(new_n291_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  OAI22_X1  g114(.A1(new_n300_), .A2(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n296_), .A2(KEYINPUT82), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318_));
  AOI21_X1  g117(.A(G176gat), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT22), .B1(new_n296_), .B2(KEYINPUT82), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n319_), .A2(new_n320_), .B1(G169gat), .B2(G176gat), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT83), .B1(new_n315_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n312_), .A2(new_n314_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT24), .B1(new_n298_), .B2(new_n291_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n278_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n309_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n316_), .A2(new_n321_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n265_), .B1(new_n323_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n255_), .B1(new_n304_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n265_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n323_), .B2(new_n330_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n303_), .A2(new_n265_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT20), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n332_), .B1(new_n336_), .B2(new_n255_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT101), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT20), .B(new_n255_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n255_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT20), .B1(new_n303_), .B2(new_n333_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n331_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n342_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n350_), .A3(KEYINPUT27), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n342_), .A3(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n352_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n253_), .B(new_n351_), .C1(new_n356_), .C2(KEYINPUT27), .ZN(new_n357_));
  INV_X1    g156(.A(new_n309_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n358_), .A2(new_n278_), .A3(new_n325_), .ZN(new_n359_));
  AOI221_X4 g158(.A(KEYINPUT83), .B1(new_n316_), .B2(new_n321_), .C1(new_n359_), .C2(new_n324_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n328_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT30), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G71gat), .B(G99gat), .ZN(new_n363_));
  INV_X1    g162(.A(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(G15gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n365_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n323_), .A2(new_n370_), .A3(new_n330_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT84), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT84), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n362_), .A2(new_n371_), .A3(new_n374_), .A4(new_n369_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n369_), .B1(new_n362_), .B2(new_n371_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT31), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT31), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n227_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n384_));
  AOI211_X1 g183(.A(KEYINPUT31), .B(new_n377_), .C1(new_n373_), .C2(new_n375_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n228_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n267_), .A2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n265_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n389_), .A2(new_n390_), .B1(new_n392_), .B2(KEYINPUT89), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(KEYINPUT89), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n217_), .A2(new_n401_), .A3(new_n223_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT28), .ZN(new_n403_));
  XOR2_X1   g202(.A(G22gat), .B(G50gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n399_), .B2(KEYINPUT91), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n397_), .B(new_n399_), .C1(KEYINPUT91), .C2(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n387_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n383_), .A2(new_n386_), .A3(new_n409_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n357_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n342_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n337_), .A2(KEYINPUT32), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n345_), .A2(new_n348_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n342_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n252_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT100), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n248_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n238_), .A2(KEYINPUT97), .A3(KEYINPUT33), .A4(new_n244_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n233_), .A2(new_n234_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n231_), .A2(new_n232_), .A3(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n237_), .A2(G225gat), .A3(G233gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n243_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n423_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT98), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n248_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT98), .B1(new_n238_), .B2(new_n244_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n422_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n354_), .A2(new_n429_), .A3(new_n355_), .A4(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT100), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n415_), .A2(new_n252_), .A3(new_n418_), .A4(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n420_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n437_), .A2(new_n387_), .A3(new_n409_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n413_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT103), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G232gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  INV_X1    g245(.A(G85gat), .ZN(new_n447_));
  INV_X1    g246(.A(G92gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n446_), .B1(new_n449_), .B2(KEYINPUT9), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT65), .B(G92gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n447_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n452_), .B2(KEYINPUT9), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT10), .B(G99gat), .Z(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT64), .B(G106gat), .Z(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT66), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n449_), .A2(new_n446_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465_));
  INV_X1    g264(.A(G99gat), .ZN(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n470_), .B2(new_n458_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT8), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT66), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n453_), .A2(new_n461_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n463_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n445_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n463_), .A2(new_n472_), .A3(new_n478_), .A4(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n443_), .A2(new_n444_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n475_), .A2(new_n479_), .B1(new_n444_), .B2(new_n443_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT71), .B1(new_n475_), .B2(new_n479_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n487_), .B(new_n483_), .C1(new_n488_), .C2(new_n445_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G190gat), .B(G218gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G134gat), .B(G162gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT36), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT72), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n486_), .A2(new_n489_), .A3(new_n496_), .A4(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n486_), .A2(new_n489_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n492_), .B(KEYINPUT36), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n439_), .A2(new_n440_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT27), .B1(new_n354_), .B2(new_n355_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n351_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n252_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n383_), .A2(new_n386_), .A3(new_n409_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n409_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n437_), .A2(new_n387_), .A3(new_n409_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT103), .B1(new_n512_), .B2(new_n502_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n504_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n515_));
  XOR2_X1   g314(.A(G71gat), .B(G78gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(KEYINPUT11), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n516_), .B(KEYINPUT67), .C1(KEYINPUT11), .C2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n475_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT12), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n523_), .A2(new_n524_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n463_), .A2(new_n474_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n472_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n475_), .A2(new_n525_), .A3(KEYINPUT12), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n531_), .A2(new_n526_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n532_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT5), .ZN(new_n538_));
  XOR2_X1   g337(.A(G176gat), .B(G204gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT68), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n536_), .A2(new_n540_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n542_), .A2(new_n543_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n515_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G1gat), .A2(G8gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT14), .ZN(new_n552_));
  INV_X1    g351(.A(G22gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G15gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n367_), .A2(G22gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n556_), .A2(KEYINPUT75), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(KEYINPUT75), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G1gat), .B(G8gat), .ZN(new_n559_));
  OR3_X1    g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n478_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT77), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(new_n561_), .A3(new_n478_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(KEYINPUT77), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n550_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n479_), .A2(new_n562_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n569_), .A2(new_n566_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n550_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n573_), .B(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n542_), .A2(new_n543_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n545_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(KEYINPUT13), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n562_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n525_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n584_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n584_), .A2(new_n590_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n549_), .A2(new_n578_), .A3(new_n581_), .A4(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n514_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G1gat), .B1(new_n599_), .B2(new_n253_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n549_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n512_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n594_), .B(KEYINPUT76), .Z(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n604_), .A2(new_n605_), .A3(KEYINPUT74), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n498_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n495_), .A2(new_n604_), .A3(new_n497_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n498_), .A2(new_n610_), .A3(new_n501_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n609_), .A2(new_n501_), .B1(new_n605_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n603_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n602_), .A2(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n615_), .A2(G1gat), .A3(new_n253_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT38), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n600_), .A2(new_n617_), .ZN(G1324gat));
  NOR2_X1   g417(.A1(new_n505_), .A2(new_n506_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n615_), .A2(G8gat), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n597_), .B(new_n621_), .C1(new_n504_), .C2(new_n513_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(KEYINPUT104), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627_));
  AOI211_X1 g426(.A(new_n627_), .B(new_n623_), .C1(new_n622_), .C2(G8gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT40), .B(new_n620_), .C1(new_n626_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1325gat));
  INV_X1    g432(.A(new_n387_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n367_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n615_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n367_), .B1(new_n598_), .B2(new_n634_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n638_), .B2(new_n637_), .ZN(G1326gat));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n598_), .A2(new_n410_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(G22gat), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT42), .B(new_n553_), .C1(new_n598_), .C2(new_n410_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n410_), .A2(new_n553_), .ZN(new_n645_));
  OAI22_X1  g444(.A1(new_n643_), .A2(new_n644_), .B1(new_n615_), .B2(new_n645_), .ZN(G1327gat));
  NOR2_X1   g445(.A1(new_n603_), .A2(new_n502_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n602_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n602_), .A2(KEYINPUT105), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n252_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n612_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(new_n612_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n512_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n603_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n601_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n663_), .A2(G29gat), .A3(new_n252_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n659_), .A2(KEYINPUT44), .A3(new_n601_), .A4(new_n660_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n654_), .B1(new_n664_), .B2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(G36gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n619_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n650_), .A2(new_n667_), .A3(new_n621_), .A4(new_n651_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT45), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(new_n672_), .A3(KEYINPUT46), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n671_), .B(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n676_), .B2(new_n669_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(new_n677_), .ZN(G1329gat));
  NAND4_X1  g477(.A1(new_n663_), .A2(G43gat), .A3(new_n634_), .A4(new_n665_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n364_), .B1(new_n652_), .B2(new_n387_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1330gat));
  OR3_X1    g482(.A1(new_n652_), .A2(G50gat), .A3(new_n409_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n663_), .A2(new_n410_), .A3(new_n665_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G50gat), .B1(new_n685_), .B2(new_n686_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1331gat));
  AND2_X1   g488(.A1(new_n549_), .A2(new_n581_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n660_), .A3(new_n578_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n514_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n253_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n690_), .A2(new_n578_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(new_n512_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n614_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n253_), .A2(G57gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1332gat));
  INV_X1    g497(.A(new_n696_), .ZN(new_n699_));
  INV_X1    g498(.A(G64gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n621_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702_));
  INV_X1    g501(.A(new_n692_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n621_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n704_), .B2(G64gat), .ZN(new_n705_));
  AOI211_X1 g504(.A(KEYINPUT48), .B(new_n700_), .C1(new_n703_), .C2(new_n621_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(G1333gat));
  OR3_X1    g506(.A1(new_n696_), .A2(G71gat), .A3(new_n387_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n634_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G71gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(G78gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n699_), .A2(new_n714_), .A3(new_n410_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n703_), .A2(new_n410_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(G78gat), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT50), .B(new_n714_), .C1(new_n703_), .C2(new_n410_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1335gat));
  NAND2_X1  g519(.A1(new_n695_), .A2(new_n647_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n447_), .B1(new_n721_), .B2(new_n253_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT108), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n656_), .B1(new_n512_), .B2(new_n657_), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT43), .B(new_n612_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n660_), .B(new_n694_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n447_), .A3(new_n253_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1336gat));
  OAI21_X1  g527(.A(new_n448_), .B1(new_n721_), .B2(new_n619_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n619_), .A2(new_n451_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n726_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT109), .Z(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n726_), .B2(new_n387_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n634_), .A2(new_n459_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n721_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(G106gat), .C1(new_n726_), .C2(new_n409_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n659_), .A2(new_n410_), .A3(new_n660_), .A4(new_n694_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT110), .A3(new_n737_), .A4(G106gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(G106gat), .B1(new_n726_), .B2(new_n409_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT52), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n695_), .A2(new_n460_), .A3(new_n410_), .A4(new_n647_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT53), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n749_), .A3(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1339gat));
  INV_X1    g550(.A(new_n578_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n549_), .A2(new_n752_), .A3(new_n581_), .ZN(new_n753_));
  OR3_X1    g552(.A1(new_n613_), .A2(KEYINPUT54), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT54), .B1(new_n613_), .B2(new_n753_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n578_), .A2(new_n546_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n475_), .A2(new_n525_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n527_), .B2(new_n526_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n759_), .A2(KEYINPUT55), .A3(new_n532_), .A4(new_n533_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n528_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(G230gat), .A3(G233gat), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n534_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n541_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n541_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT111), .B(KEYINPUT56), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n766_), .A2(KEYINPUT112), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(KEYINPUT112), .A3(new_n768_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n757_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n565_), .A2(new_n550_), .A3(new_n567_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n570_), .A2(new_n571_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n576_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT113), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n577_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n773_), .A2(new_n774_), .A3(new_n778_), .A4(new_n576_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n502_), .B1(new_n772_), .B2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n780_), .A2(new_n545_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n766_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n541_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n612_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n785_), .B(KEYINPUT58), .C1(new_n786_), .C2(new_n787_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n782_), .A2(new_n783_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT57), .B(new_n502_), .C1(new_n772_), .C2(new_n781_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n771_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n578_), .B(new_n546_), .C1(new_n769_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n781_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n503_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT115), .B1(new_n798_), .B2(KEYINPUT57), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n791_), .B1(new_n794_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n594_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n756_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n619_), .A2(new_n252_), .ZN(new_n803_));
  OR3_X1    g602(.A1(new_n803_), .A2(KEYINPUT116), .A3(new_n412_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n803_), .B2(new_n412_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n802_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n578_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n754_), .A2(new_n755_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n788_), .A2(new_n784_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n657_), .A2(new_n811_), .A3(new_n790_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n783_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n798_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n792_), .A2(new_n793_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n798_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n810_), .B1(new_n817_), .B2(new_n594_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n806_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n809_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n756_), .B1(new_n800_), .B2(new_n660_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n819_), .A2(KEYINPUT117), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n819_), .A2(KEYINPUT117), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n809_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n578_), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT118), .B2(G113gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n808_), .B1(new_n826_), .B2(new_n828_), .ZN(G1340gat));
  INV_X1    g628(.A(new_n690_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n818_), .A2(new_n819_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n820_), .A2(new_n825_), .A3(new_n690_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n832_), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n807_), .A2(new_n840_), .A3(new_n603_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n820_), .A2(new_n825_), .A3(new_n801_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n840_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n818_), .A2(new_n819_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n502_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n821_), .A2(new_n824_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n612_), .A2(new_n844_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n849_), .B(new_n850_), .C1(new_n807_), .C2(new_n809_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT120), .B(new_n844_), .C1(new_n845_), .C2(new_n502_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n848_), .A2(new_n851_), .A3(new_n852_), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n803_), .A2(new_n411_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT121), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n802_), .A2(KEYINPUT122), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  INV_X1    g656(.A(new_n855_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n818_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n578_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G141gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT122), .B1(new_n802_), .B2(new_n855_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n818_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(G141gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n578_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(G1344gat));
  OAI21_X1  g666(.A(new_n830_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G148gat), .ZN(new_n869_));
  INV_X1    g668(.A(G148gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n870_), .A3(new_n830_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1345gat));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT123), .Z(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n864_), .B2(new_n603_), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n660_), .B(new_n874_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1346gat));
  NAND3_X1  g677(.A1(new_n864_), .A2(new_n203_), .A3(new_n503_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n612_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n203_), .B2(new_n880_), .ZN(G1347gat));
  OAI21_X1  g680(.A(new_n810_), .B1(new_n817_), .B2(new_n603_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n621_), .A2(new_n253_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(new_n387_), .A3(new_n410_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885_), .B2(new_n752_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT62), .B(G169gat), .C1(new_n885_), .C2(new_n752_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n885_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n578_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n888_), .B(new_n889_), .C1(new_n269_), .C2(new_n891_), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n890_), .B2(new_n830_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n802_), .A2(new_n410_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n690_), .A2(new_n883_), .A3(new_n297_), .A4(new_n387_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(new_n898_), .A3(new_n895_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n893_), .B1(new_n897_), .B2(new_n899_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n660_), .A2(new_n387_), .A3(new_n883_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G183gat), .B1(new_n894_), .B2(new_n901_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n594_), .A2(new_n288_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n890_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n885_), .B2(new_n612_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n502_), .A2(new_n283_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n885_), .B2(new_n906_), .ZN(G1351gat));
  NOR3_X1   g706(.A1(new_n802_), .A2(new_n411_), .A3(new_n883_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n578_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n830_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT125), .B(G204gat), .Z(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n908_), .A2(KEYINPUT125), .A3(G204gat), .A4(new_n830_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1353gat));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n916_));
  INV_X1    g715(.A(G211gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n594_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT126), .Z(new_n919_));
  NAND2_X1  g718(.A1(new_n908_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n916_), .A2(new_n917_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1354gat));
  NAND2_X1  g721(.A1(new_n908_), .A2(new_n503_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT127), .B(G218gat), .Z(new_n924_));
  NOR2_X1   g723(.A1(new_n612_), .A2(new_n924_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n923_), .A2(new_n924_), .B1(new_n908_), .B2(new_n925_), .ZN(G1355gat));
endmodule


