//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT6), .Z(new_n209_));
  XNOR2_X1  g008(.A(G85gat), .B(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NOR4_X1   g014(.A1(new_n207_), .A2(new_n209_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n217_), .B2(KEYINPUT8), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n209_), .B2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n217_), .A2(KEYINPUT8), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n223_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n216_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G29gat), .B(G36gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT15), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  AOI211_X1 g031(.A(new_n204_), .B(new_n232_), .C1(new_n229_), .C2(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  XOR2_X1   g034(.A(G190gat), .B(G218gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT70), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G134gat), .B(G162gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n240_), .A2(KEYINPUT36), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT71), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT72), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n233_), .B(new_n234_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(KEYINPUT36), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT37), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n244_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(new_n246_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT73), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G57gat), .B(G64gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT11), .ZN(new_n257_));
  XOR2_X1   g056(.A(G71gat), .B(G78gat), .Z(new_n258_));
  OR2_X1    g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n256_), .A2(KEYINPUT11), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G231gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G8gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G15gat), .ZN(new_n268_));
  INV_X1    g067(.A(G22gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G15gat), .A2(G22gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G1gat), .A2(G8gat), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n270_), .A2(new_n271_), .B1(KEYINPUT14), .B2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n267_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n267_), .A2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n264_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT75), .ZN(new_n278_));
  XOR2_X1   g077(.A(G127gat), .B(G155gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT16), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G183gat), .B(G211gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT17), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT76), .Z(new_n285_));
  INV_X1    g084(.A(KEYINPUT17), .ZN(new_n286_));
  OR3_X1    g085(.A1(new_n277_), .A2(new_n286_), .A3(new_n282_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n255_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT64), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n226_), .A2(new_n262_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n226_), .A2(new_n262_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT66), .ZN(new_n297_));
  INV_X1    g096(.A(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n295_), .B1(new_n304_), .B2(new_n302_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n297_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT5), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n297_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(KEYINPUT13), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n290_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n276_), .A2(new_n230_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n267_), .B(new_n273_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n229_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G229gat), .A2(G233gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT78), .Z(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT77), .B1(new_n325_), .B2(new_n229_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n325_), .A2(new_n229_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G229gat), .A3(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G113gat), .B(G141gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G169gat), .B(G197gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(G78gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(new_n206_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT88), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n348_), .A2(KEYINPUT1), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(KEYINPUT1), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(G141gat), .ZN(new_n354_));
  INV_X1    g153(.A(G148gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n352_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n348_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(new_n351_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT3), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n359_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT87), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n360_), .A2(new_n362_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT86), .B1(new_n372_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n359_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n357_), .B1(new_n371_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n347_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n347_), .A3(new_n383_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n346_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n388_), .A2(KEYINPUT88), .A3(new_n384_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n345_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT88), .B1(new_n388_), .B2(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n385_), .A2(new_n346_), .A3(new_n386_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n345_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT90), .B(G197gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G204gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n398_));
  INV_X1    g197(.A(G204gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n401_));
  INV_X1    g200(.A(G197gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(G204gat), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n397_), .A2(new_n398_), .A3(new_n400_), .A4(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G211gat), .B(G218gat), .Z(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n399_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT21), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(G197gat), .B2(G204gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n397_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n405_), .A2(KEYINPUT21), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n404_), .A2(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT89), .ZN(new_n415_));
  XOR2_X1   g214(.A(G22gat), .B(G50gat), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n414_), .A2(KEYINPUT89), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(KEYINPUT89), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n395_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n390_), .A2(new_n417_), .A3(new_n421_), .A4(new_n394_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT82), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT22), .B(G169gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT23), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(G183gat), .A3(G190gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G183gat), .A2(G190gat), .ZN(new_n434_));
  OAI221_X1 g233(.A(new_n427_), .B1(new_n428_), .B2(G176gat), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(KEYINPUT83), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n429_), .A2(new_n437_), .A3(KEYINPUT23), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n432_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT80), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT26), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n441_), .A2(new_n442_), .A3(G190gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G190gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G183gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT25), .B1(new_n446_), .B2(KEYINPUT79), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n446_), .A2(KEYINPUT25), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(KEYINPUT79), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n440_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G169gat), .A2(G176gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT24), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n427_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(KEYINPUT24), .A3(new_n454_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n435_), .B1(new_n450_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G43gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n461_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G127gat), .B(G134gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G113gat), .B(G120gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT84), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT85), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n464_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(new_n268_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT30), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT31), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n471_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n425_), .A2(new_n477_), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n382_), .A2(KEYINPUT4), .A3(new_n469_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G225gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n382_), .B2(new_n469_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n357_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n380_), .B1(new_n379_), .B2(new_n359_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n359_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT87), .B(new_n488_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n469_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(KEYINPUT95), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n468_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n465_), .A2(new_n466_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n496_), .B(new_n357_), .C1(new_n371_), .C2(new_n381_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AND4_X1   g297(.A1(KEYINPUT96), .A2(new_n493_), .A3(KEYINPUT4), .A4(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n485_), .B2(new_n492_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT96), .B1(new_n500_), .B2(KEYINPUT4), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n483_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n480_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT97), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT97), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n505_), .A3(new_n480_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G29gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G85gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT0), .B(G57gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  NAND4_X1  g310(.A1(new_n502_), .A2(new_n507_), .A3(KEYINPUT33), .A4(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n461_), .B2(new_n413_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G226gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT19), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n428_), .A2(KEYINPUT94), .ZN(new_n518_));
  INV_X1    g317(.A(G176gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT22), .B(G169gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n519_), .A3(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n446_), .A2(KEYINPUT23), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n436_), .A2(new_n438_), .B1(G190gat), .B2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n523_), .B(new_n427_), .C1(new_n434_), .C2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n444_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT25), .B(G183gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n444_), .A2(new_n527_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n453_), .A2(KEYINPUT24), .A3(new_n426_), .A4(new_n454_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n433_), .B1(new_n456_), .B2(new_n451_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n514_), .B(new_n517_), .C1(new_n413_), .C2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT20), .B1(new_n461_), .B2(new_n413_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n412_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n516_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G8gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT18), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G64gat), .B(G92gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n536_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n480_), .B(new_n479_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n511_), .B1(new_n500_), .B2(new_n481_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n493_), .A2(KEYINPUT4), .A3(new_n498_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n500_), .A2(KEYINPUT96), .A3(KEYINPUT4), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n482_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AND4_X1   g355(.A1(new_n505_), .A2(new_n493_), .A3(new_n498_), .A4(new_n480_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n505_), .B1(new_n500_), .B2(new_n480_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n511_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n556_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n512_), .B(new_n551_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT99), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n535_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n526_), .A2(new_n534_), .A3(KEYINPUT99), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n412_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n517_), .B1(new_n568_), .B2(new_n514_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n537_), .A2(new_n516_), .A3(new_n538_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n544_), .A2(KEYINPUT32), .ZN(new_n572_));
  MUX2_X1   g371(.A(new_n571_), .B(new_n540_), .S(new_n572_), .Z(new_n573_));
  AOI21_X1  g372(.A(new_n511_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n561_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n478_), .B1(new_n564_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n547_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n545_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n547_), .A2(new_n577_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT27), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n548_), .A2(KEYINPUT27), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n560_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n502_), .A2(new_n511_), .A3(new_n507_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n423_), .A2(new_n477_), .A3(new_n424_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n424_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n390_), .A2(new_n394_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n476_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n576_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n323_), .A2(new_n341_), .A3(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n561_), .A2(new_n574_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n594_), .A2(G1gat), .A3(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT38), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n244_), .A2(new_n247_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n593_), .A2(new_n289_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n341_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n322_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n603_), .B2(new_n595_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n598_), .A3(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(G8gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n603_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n584_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT39), .A3(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n594_), .A2(G8gat), .A3(new_n584_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(G1325gat));
  OAI21_X1  g418(.A(G15gat), .B1(new_n603_), .B2(new_n477_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT41), .Z(new_n621_));
  INV_X1    g420(.A(new_n594_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n268_), .A3(new_n476_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1326gat));
  OAI21_X1  g423(.A(G22gat), .B1(new_n603_), .B2(new_n425_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n425_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n622_), .A2(new_n269_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n599_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n288_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n322_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n593_), .A3(new_n341_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(G29gat), .A3(new_n595_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n254_), .B1(new_n576_), .B2(new_n592_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n254_), .B(KEYINPUT43), .C1(new_n576_), .C2(new_n592_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(new_n288_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT44), .A4(new_n602_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n638_), .A2(new_n288_), .A3(new_n602_), .A4(new_n639_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT104), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT44), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n289_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(KEYINPUT103), .A3(new_n602_), .A4(new_n639_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n642_), .A2(new_n645_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n595_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n635_), .B1(new_n652_), .B2(G29gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT105), .ZN(G1328gat));
  NOR3_X1   g453(.A1(new_n634_), .A2(G36gat), .A3(new_n584_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT45), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n642_), .A2(new_n645_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n643_), .A2(new_n646_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n608_), .A4(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n658_), .B1(new_n650_), .B2(new_n608_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n656_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT107), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(KEYINPUT107), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n657_), .A2(new_n608_), .A3(new_n660_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(G36gat), .A3(new_n661_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n671_), .A2(KEYINPUT107), .A3(new_n665_), .A4(new_n656_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n668_), .A2(new_n672_), .ZN(G1329gat));
  NAND3_X1  g472(.A1(new_n650_), .A2(G43gat), .A3(new_n476_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n634_), .A2(new_n477_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(G43gat), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n676_), .B(new_n677_), .Z(G1330gat));
  INV_X1    g477(.A(G50gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n628_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT110), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n634_), .A2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT109), .B(new_n679_), .C1(new_n650_), .C2(new_n628_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n657_), .A2(new_n628_), .A3(new_n660_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(G50gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT111), .B(new_n682_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n321_), .A2(new_n341_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n600_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G57gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n595_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n593_), .A2(new_n601_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n696_), .A2(new_n322_), .A3(new_n289_), .A4(new_n255_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT112), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT112), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n651_), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n695_), .B1(new_n701_), .B2(new_n694_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n703_), .A3(new_n608_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n693_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n705_), .B2(new_n608_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n706_), .A2(new_n707_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n704_), .B1(new_n709_), .B2(new_n710_), .ZN(G1333gat));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n698_), .A2(new_n712_), .A3(new_n476_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n705_), .B2(new_n476_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n714_), .A2(new_n715_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(G1334gat));
  NAND3_X1  g518(.A1(new_n698_), .A2(new_n343_), .A3(new_n628_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n343_), .B1(new_n705_), .B2(new_n628_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n721_), .A2(new_n722_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n724_), .B2(new_n725_), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n640_), .A2(new_n692_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n595_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n632_), .A2(new_n321_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n696_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(new_n213_), .A3(new_n651_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1336gat));
  OAI21_X1  g532(.A(G92gat), .B1(new_n727_), .B2(new_n584_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n214_), .A3(new_n608_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT115), .Z(G1337gat));
  OAI21_X1  g536(.A(G99gat), .B1(new_n727_), .B2(new_n477_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n731_), .A2(new_n476_), .A3(new_n205_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n740_), .B(new_n741_), .Z(G1338gat));
  NOR3_X1   g541(.A1(new_n730_), .A2(G106gat), .A3(new_n425_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT117), .Z(new_n744_));
  OAI21_X1  g543(.A(G106gat), .B1(new_n727_), .B2(new_n425_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g549(.A(G113gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n307_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n303_), .A2(new_n305_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n292_), .B1(new_n754_), .B2(new_n294_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n301_), .A2(new_n306_), .A3(KEYINPUT55), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n312_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n312_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n332_), .A2(new_n327_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n324_), .A2(new_n326_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n762_), .B(new_n338_), .C1(new_n327_), .C2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n340_), .A2(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(KEYINPUT120), .A3(new_n315_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT120), .B1(new_n765_), .B2(new_n315_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n760_), .A2(new_n761_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n760_), .B2(new_n768_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n254_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n757_), .A2(new_n312_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n312_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n341_), .A2(new_n315_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n759_), .B2(KEYINPUT118), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n780_), .A2(KEYINPUT119), .B1(new_n316_), .B2(new_n765_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n777_), .A2(new_n782_), .A3(new_n779_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n631_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n771_), .B1(new_n784_), .B2(KEYINPUT57), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n786_), .B(new_n631_), .C1(new_n781_), .C2(new_n783_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n288_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n323_), .A2(new_n601_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT54), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n591_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n595_), .A2(new_n608_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n751_), .B1(new_n794_), .B2(new_n601_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT121), .B(new_n751_), .C1(new_n794_), .C2(new_n601_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n591_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT59), .A3(new_n793_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n601_), .A2(new_n751_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n797_), .A2(new_n798_), .B1(new_n803_), .B2(new_n804_), .ZN(G1340gat));
  INV_X1    g604(.A(new_n794_), .ZN(new_n806_));
  XOR2_X1   g605(.A(KEYINPUT122), .B(G120gat), .Z(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n321_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n806_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n807_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n321_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n807_), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n812_), .A3(new_n289_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n288_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n812_), .ZN(G1342gat));
  INV_X1    g614(.A(G134gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n794_), .B2(new_n599_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT123), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n816_), .C1(new_n794_), .C2(new_n599_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n255_), .A2(new_n816_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n818_), .A2(new_n820_), .B1(new_n803_), .B2(new_n821_), .ZN(G1343gat));
  INV_X1    g621(.A(new_n588_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n769_), .A2(new_n254_), .A3(new_n770_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT118), .ZN(new_n825_));
  INV_X1    g624(.A(new_n778_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n316_), .A2(new_n765_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n783_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n599_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n824_), .B1(new_n831_), .B2(new_n786_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n784_), .A2(KEYINPUT57), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n289_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n789_), .B(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n823_), .B(new_n793_), .C1(new_n834_), .C2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n601_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(new_n354_), .ZN(G1344gat));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n321_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(new_n355_), .ZN(G1345gat));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n288_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n842_), .B(new_n843_), .Z(G1346gat));
  OAI21_X1  g643(.A(G162gat), .B1(new_n837_), .B2(new_n255_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n588_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n599_), .A2(G162gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n793_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n845_), .A2(KEYINPUT124), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1347gat));
  NOR2_X1   g652(.A1(new_n651_), .A2(new_n584_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n792_), .B(new_n854_), .C1(new_n834_), .C2(new_n836_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G169gat), .B1(new_n855_), .B2(new_n601_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n791_), .A2(new_n341_), .A3(new_n792_), .A4(new_n854_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(KEYINPUT125), .A3(G169gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(KEYINPUT62), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n518_), .A2(new_n522_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT125), .B1(new_n859_), .B2(G169gat), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(G1348gat));
  NOR2_X1   g666(.A1(new_n855_), .A2(new_n321_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n519_), .A2(KEYINPUT126), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n519_), .A2(KEYINPUT126), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n868_), .B2(new_n870_), .ZN(G1349gat));
  NOR2_X1   g671(.A1(new_n855_), .A2(new_n288_), .ZN(new_n873_));
  MUX2_X1   g672(.A(G183gat), .B(new_n529_), .S(new_n873_), .Z(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n855_), .B2(new_n255_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n631_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n855_), .B2(new_n876_), .ZN(G1351gat));
  NAND2_X1  g676(.A1(new_n846_), .A2(new_n854_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n601_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n402_), .ZN(G1352gat));
  INV_X1    g679(.A(new_n878_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n322_), .C1(KEYINPUT127), .C2(new_n399_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT127), .B(G204gat), .Z(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n878_), .B2(new_n321_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1353gat));
  XOR2_X1   g684(.A(KEYINPUT63), .B(G211gat), .Z(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(new_n289_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n878_), .B2(new_n288_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1354gat));
  OAI21_X1  g689(.A(G218gat), .B1(new_n878_), .B2(new_n255_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n599_), .A2(G218gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n878_), .B2(new_n892_), .ZN(G1355gat));
endmodule


