//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OR2_X1    g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT94), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G211gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G218gat), .ZN(new_n210_));
  INV_X1    g009(.A(G218gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(G211gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT95), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(G211gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(G218gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT95), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n204_), .A2(new_n205_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n208_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT96), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n216_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n213_), .A2(KEYINPUT96), .A3(new_n217_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n206_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT97), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT97), .A4(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n223_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G141gat), .A2(G148gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(KEYINPUT1), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G155gat), .A3(G162gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n249_), .A3(new_n244_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G141gat), .B(G148gat), .Z(new_n251_));
  AOI22_X1  g050(.A1(new_n243_), .A2(new_n246_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n203_), .B1(new_n234_), .B2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n208_), .A2(new_n222_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n206_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT97), .B1(new_n257_), .B2(new_n228_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n233_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n256_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n243_), .A2(new_n246_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n250_), .A2(new_n251_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT29), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT93), .B1(new_n252_), .B2(new_n253_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n202_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n255_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT98), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT28), .B1(new_n263_), .B2(KEYINPUT29), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n252_), .A2(new_n274_), .A3(new_n253_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G22gat), .B(G50gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n276_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n270_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n255_), .A2(new_n268_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT99), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT98), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n269_), .A2(new_n284_), .A3(new_n270_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n255_), .A2(new_n268_), .A3(KEYINPUT99), .A4(new_n280_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n272_), .A2(new_n283_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n271_), .A2(new_n281_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n279_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT100), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT22), .B(G169gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT88), .B(G176gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(G183gat), .B2(G190gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(G183gat), .A3(G190gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT86), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n300_), .A2(new_n296_), .A3(G183gat), .A4(G190gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n297_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n292_), .B(new_n295_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G183gat), .ZN(new_n308_));
  INV_X1    g107(.A(G190gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT23), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n298_), .ZN(new_n311_));
  INV_X1    g110(.A(G169gat), .ZN(new_n312_));
  INV_X1    g111(.A(G176gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT24), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n307_), .A2(new_n311_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n304_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(new_n256_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT20), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT19), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n307_), .A2(new_n316_), .A3(new_n315_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(new_n302_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(G169gat), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n294_), .B(new_n328_), .C1(new_n293_), .C2(new_n326_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n292_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  INV_X1    g130(.A(new_n303_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n311_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n311_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n325_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n323_), .B1(new_n234_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n291_), .B1(new_n320_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT20), .B1(new_n234_), .B2(new_n318_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n232_), .A2(new_n233_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n340_), .A2(new_n256_), .A3(new_n336_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n322_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n234_), .B2(new_n318_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n336_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n260_), .A2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n344_), .A2(new_n346_), .A3(KEYINPUT100), .A4(new_n323_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n338_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n338_), .A2(new_n342_), .A3(new_n347_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n339_), .A2(new_n341_), .A3(new_n322_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n323_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n352_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT104), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n234_), .A2(new_n336_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n322_), .B1(new_n320_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n318_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n260_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n234_), .A2(new_n336_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT20), .A4(new_n323_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n354_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT104), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n362_), .A2(KEYINPUT27), .A3(new_n371_), .A4(new_n355_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G71gat), .B(G99gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G43gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT92), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n381_));
  INV_X1    g180(.A(new_n377_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n378_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n377_), .A2(new_n378_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n380_), .A2(new_n381_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n381_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n377_), .A2(new_n378_), .A3(new_n385_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n376_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT31), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n336_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n336_), .A2(new_n399_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n395_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n404_), .A2(KEYINPUT31), .A3(new_n400_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n394_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT31), .B1(new_n404_), .B2(new_n400_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n393_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n392_), .A2(new_n263_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n252_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n263_), .B1(new_n384_), .B2(new_n379_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT4), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n414_), .A2(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n417_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G85gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT0), .B(G57gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n419_), .A2(new_n421_), .A3(KEYINPUT103), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(new_n421_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT103), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n419_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n410_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  AND4_X1   g232(.A1(new_n290_), .A2(new_n358_), .A3(new_n372_), .A4(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n338_), .A2(new_n342_), .A3(new_n347_), .A4(new_n435_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n432_), .A2(new_n437_), .A3(new_n438_), .A4(new_n427_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n420_), .A2(new_n417_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n425_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT102), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n413_), .A2(new_n416_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(new_n417_), .ZN(new_n444_));
  AOI211_X1 g243(.A(KEYINPUT102), .B(new_n418_), .C1(new_n413_), .C2(new_n416_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n441_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n428_), .A2(new_n425_), .B1(KEYINPUT101), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(KEYINPUT101), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n426_), .B(new_n449_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n439_), .B1(new_n356_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n290_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n287_), .A2(new_n289_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n358_), .A3(new_n372_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n434_), .B1(new_n456_), .B2(new_n410_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G113gat), .B(G141gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G169gat), .B(G197gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G8gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n470_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n466_), .B(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n472_), .A3(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n480_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n473_), .B(new_n484_), .Z(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n485_), .B2(new_n468_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n473_), .B(new_n484_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(KEYINPUT84), .A3(new_n475_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n482_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n461_), .B1(new_n481_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n477_), .B(KEYINPUT83), .ZN(new_n492_));
  INV_X1    g291(.A(new_n480_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n494_), .A3(new_n460_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n496_), .B(KEYINPUT85), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n457_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G230gat), .A2(G233gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT64), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n503_));
  INV_X1    g302(.A(G85gat), .ZN(new_n504_));
  INV_X1    g303(.A(G92gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT10), .B(G99gat), .Z(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT66), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n508_), .A2(new_n509_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n514_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT67), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n526_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n534_), .A3(new_n519_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n506_), .A2(new_n507_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT8), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n521_), .A2(new_n532_), .A3(new_n526_), .A4(new_n522_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n536_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n525_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G78gat), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n502_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n538_), .A2(new_n541_), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n514_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n542_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n550_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n560_), .B(new_n550_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n552_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT68), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n554_), .A2(new_n555_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n562_), .A2(new_n563_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n502_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n561_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT70), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT72), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n569_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT37), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT36), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT76), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT34), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(KEYINPUT35), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n542_), .B2(new_n473_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n542_), .A2(new_n485_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(KEYINPUT74), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n554_), .A2(new_n487_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n591_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n600_));
  INV_X1    g399(.A(new_n591_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n542_), .B2(new_n485_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n541_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n540_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n553_), .B(new_n473_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n592_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n600_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n593_), .A2(new_n596_), .A3(KEYINPUT75), .A4(new_n601_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n586_), .B1(new_n599_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n599_), .A2(new_n610_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n581_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n599_), .A2(new_n610_), .A3(new_n613_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n585_), .B1(new_n599_), .B2(new_n610_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n616_), .A2(new_n617_), .A3(KEYINPUT37), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT77), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n610_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n607_), .B1(new_n597_), .B2(new_n596_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n594_), .A2(KEYINPUT74), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n601_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n581_), .B(new_n614_), .C1(new_n624_), .C2(new_n585_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n611_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT77), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n619_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n475_), .B(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(new_n555_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n555_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT78), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT78), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n636_), .A2(new_n638_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n643_), .B(KEYINPUT17), .Z(new_n646_));
  NAND2_X1  g445(.A1(new_n635_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT81), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n635_), .A2(KEYINPUT81), .A3(new_n646_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT82), .Z(new_n652_));
  NOR3_X1   g451(.A1(new_n580_), .A2(new_n629_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n499_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT105), .Z(new_n655_));
  NAND2_X1  g454(.A1(new_n432_), .A2(new_n427_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n463_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n616_), .A2(new_n617_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n457_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n496_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n580_), .A2(new_n663_), .A3(new_n651_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n656_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n659_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n660_), .A2(new_n666_), .A3(new_n667_), .ZN(G1324gat));
  XNOR2_X1  g467(.A(new_n369_), .B(KEYINPUT104), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n355_), .A2(KEYINPUT27), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n669_), .A2(new_n670_), .B1(new_n357_), .B2(new_n356_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n655_), .A2(new_n464_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G8gat), .B1(new_n665_), .B2(new_n671_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT39), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(KEYINPUT40), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  OAI21_X1  g479(.A(G15gat), .B1(new_n665_), .B2(new_n410_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT41), .Z(new_n682_));
  INV_X1    g481(.A(new_n410_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n397_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n654_), .B2(new_n684_), .ZN(G1326gat));
  OAI21_X1  g484(.A(G22gat), .B1(new_n665_), .B2(new_n290_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT42), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n290_), .A2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n654_), .B2(new_n688_), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n652_), .A2(new_n661_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n580_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n499_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n657_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n578_), .B(KEYINPUT13), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n496_), .A3(new_n652_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n619_), .A2(new_n628_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n683_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n629_), .B(new_n699_), .C1(new_n700_), .C2(new_n434_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(KEYINPUT44), .ZN(new_n703_));
  INV_X1    g502(.A(new_n696_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n434_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n671_), .A2(new_n454_), .B1(new_n452_), .B2(new_n290_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n683_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n699_), .B1(new_n707_), .B2(new_n629_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n701_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n704_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT106), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n702_), .A2(new_n712_), .A3(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n703_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n657_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n694_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  XNOR2_X1  g515(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n671_), .A2(G36gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n693_), .A2(KEYINPUT45), .A3(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721_));
  INV_X1    g520(.A(new_n719_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n692_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n704_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n671_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n698_), .A2(new_n701_), .ZN(new_n728_));
  AND4_X1   g527(.A1(new_n712_), .A2(new_n728_), .A3(KEYINPUT44), .A4(new_n704_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n712_), .B1(new_n702_), .B2(KEYINPUT44), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n731_), .B2(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n718_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G36gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n711_), .A2(new_n713_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n727_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT107), .B(new_n717_), .C1(new_n737_), .C2(new_n724_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n734_), .A2(new_n738_), .ZN(G1329gat));
  INV_X1    g538(.A(G43gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n410_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n714_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n692_), .B2(new_n410_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1330gat));
  INV_X1    g546(.A(G50gat), .ZN(new_n748_));
  INV_X1    g547(.A(new_n290_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n714_), .B2(new_n749_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n692_), .A2(G50gat), .A3(new_n290_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT110), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753_));
  INV_X1    g552(.A(new_n751_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n290_), .B(new_n703_), .C1(new_n711_), .C2(new_n713_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n753_), .B(new_n754_), .C1(new_n755_), .C2(new_n748_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n752_), .A2(new_n756_), .ZN(G1331gat));
  XNOR2_X1  g556(.A(new_n651_), .B(KEYINPUT82), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n697_), .A2(new_n758_), .ZN(new_n759_));
  NOR4_X1   g558(.A1(new_n759_), .A2(new_n457_), .A3(new_n496_), .A4(new_n695_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n657_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT111), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n695_), .A2(new_n652_), .A3(new_n497_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n662_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G57gat), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n656_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n762_), .A2(new_n766_), .ZN(G1332gat));
  OAI21_X1  g566(.A(G64gat), .B1(new_n764_), .B2(new_n671_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(G64gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n771_), .A3(new_n672_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n764_), .B2(new_n410_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n760_), .A2(new_n776_), .A3(new_n683_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1334gat));
  OAI21_X1  g577(.A(G78gat), .B1(new_n764_), .B2(new_n290_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT50), .ZN(new_n780_));
  INV_X1    g579(.A(G78gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n760_), .A2(new_n781_), .A3(new_n749_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n695_), .A2(new_n496_), .A3(new_n758_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n728_), .A2(KEYINPUT113), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n728_), .A2(KEYINPUT113), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787_), .B2(new_n656_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n690_), .A2(new_n695_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n707_), .A3(new_n663_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n504_), .A3(new_n657_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n792_), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n787_), .A2(new_n505_), .A3(new_n671_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n505_), .B1(new_n790_), .B2(new_n671_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT114), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n787_), .B2(new_n410_), .ZN(new_n798_));
  OR2_X1    g597(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n683_), .A2(new_n511_), .ZN(new_n801_));
  OR3_X1    g600(.A1(new_n790_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n790_), .B2(new_n801_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n802_), .A2(new_n803_), .B1(KEYINPUT116), .B2(KEYINPUT51), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n798_), .A2(new_n799_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n799_), .B1(new_n798_), .B2(new_n804_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n791_), .A2(new_n512_), .A3(new_n749_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n784_), .A2(new_n749_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n512_), .B1(new_n810_), .B2(new_n728_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n812_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n808_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g615(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n697_), .A2(new_n695_), .A3(new_n758_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n497_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n653_), .A2(new_n498_), .A3(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n559_), .A2(new_n561_), .A3(new_n568_), .A4(new_n575_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n496_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n550_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n556_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n554_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n562_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n828_), .A2(KEYINPUT55), .B1(new_n829_), .B2(new_n502_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n559_), .A2(new_n831_), .A3(new_n561_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n575_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n824_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n834_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT119), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n833_), .A2(new_n834_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n839_), .A2(new_n836_), .A3(new_n840_), .A4(new_n824_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n486_), .A2(new_n488_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n493_), .A3(new_n474_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n461_), .C1(new_n493_), .C2(new_n479_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(new_n495_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n578_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n838_), .A2(new_n841_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n661_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(KEYINPUT57), .A3(new_n848_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n833_), .B2(KEYINPUT56), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(KEYINPUT56), .B2(new_n833_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n845_), .A2(new_n823_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n833_), .A2(KEYINPUT56), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n853_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT58), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(new_n858_), .A3(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n629_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n851_), .A2(new_n852_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n822_), .B1(new_n863_), .B2(new_n651_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n671_), .A2(new_n657_), .A3(new_n290_), .A4(new_n683_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(G113gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n496_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT59), .B1(new_n864_), .B2(new_n865_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n865_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n871_), .B2(new_n865_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n861_), .A2(new_n629_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n859_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n847_), .B2(new_n848_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n758_), .B1(new_n877_), .B2(new_n852_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n878_), .B2(new_n822_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n869_), .A2(new_n497_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n868_), .B1(new_n880_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n695_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n866_), .B(new_n883_), .C1(KEYINPUT60), .C2(new_n882_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n869_), .A2(new_n580_), .A3(new_n879_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n882_), .ZN(G1341gat));
  INV_X1    g685(.A(G127gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n866_), .A2(new_n887_), .A3(new_n758_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n651_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n869_), .A2(new_n889_), .A3(new_n879_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(new_n887_), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n866_), .A2(new_n892_), .A3(new_n661_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n869_), .A2(new_n629_), .A3(new_n879_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n892_), .ZN(G1343gat));
  NOR4_X1   g694(.A1(new_n672_), .A2(new_n683_), .A3(new_n290_), .A4(new_n656_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT122), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n864_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n496_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n580_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n758_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n864_), .A2(new_n848_), .A3(new_n898_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(G162gat), .ZN(new_n909_));
  INV_X1    g708(.A(new_n822_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n847_), .A2(KEYINPUT57), .A3(new_n848_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n911_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(new_n889_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n661_), .A3(new_n897_), .ZN(new_n914_));
  INV_X1    g713(.A(G162gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(KEYINPUT123), .A3(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n697_), .A2(new_n915_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n909_), .A2(new_n916_), .B1(new_n899_), .B2(new_n917_), .ZN(G1347gat));
  AOI21_X1  g717(.A(new_n822_), .B1(new_n863_), .B2(new_n652_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n672_), .A2(new_n433_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n749_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n919_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n496_), .ZN(new_n924_));
  XOR2_X1   g723(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(G169gat), .A3(new_n926_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n919_), .A2(new_n663_), .A3(new_n922_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n925_), .B1(new_n928_), .B2(new_n312_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n293_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n929_), .A3(new_n930_), .ZN(G1348gat));
  NOR3_X1   g730(.A1(new_n919_), .A2(new_n695_), .A3(new_n922_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n294_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT125), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n580_), .B(new_n921_), .C1(new_n878_), .C2(new_n822_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n935_), .A2(new_n936_), .A3(new_n294_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n913_), .A2(new_n938_), .A3(new_n290_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT126), .B1(new_n864_), .B2(new_n749_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n695_), .A2(new_n920_), .A3(new_n313_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n934_), .A2(new_n937_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  NOR4_X1   g742(.A1(new_n919_), .A2(new_n305_), .A3(new_n651_), .A4(new_n922_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n920_), .A2(new_n652_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n938_), .B1(new_n913_), .B2(new_n290_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n864_), .A2(KEYINPUT126), .A3(new_n749_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n944_), .B1(new_n948_), .B2(new_n308_), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n923_), .A2(new_n306_), .A3(new_n661_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n919_), .A2(new_n697_), .A3(new_n922_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n309_), .ZN(G1351gat));
  NAND3_X1  g751(.A1(new_n672_), .A2(new_n454_), .A3(new_n410_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n864_), .A2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n496_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n580_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g757(.A(KEYINPUT63), .B(G211gat), .C1(new_n954_), .C2(new_n889_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(KEYINPUT63), .B(G211gat), .ZN(new_n960_));
  NOR4_X1   g759(.A1(new_n864_), .A2(new_n651_), .A3(new_n953_), .A4(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1354gat));
  AOI21_X1  g761(.A(G218gat), .B1(new_n954_), .B2(new_n661_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n629_), .A2(G218gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(KEYINPUT127), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n954_), .B2(new_n965_), .ZN(G1355gat));
endmodule


