//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n204_), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G71gat), .B(G78gat), .Z(new_n219_));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(KEYINPUT11), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT11), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n220_), .B2(KEYINPUT11), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n214_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n228_), .B(new_n216_), .C1(new_n208_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT64), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n231_), .A2(new_n232_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n228_), .B1(new_n241_), .B2(new_n216_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n234_), .B1(new_n242_), .B2(KEYINPUT65), .ZN(new_n243_));
  INV_X1    g042(.A(new_n216_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT64), .B1(new_n237_), .B2(new_n238_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(new_n233_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n246_), .B2(new_n239_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n228_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n218_), .B(new_n227_), .C1(new_n243_), .C2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n248_), .B1(new_n247_), .B2(new_n228_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n241_), .A2(new_n216_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n254_), .A3(new_n234_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n227_), .B1(new_n255_), .B2(new_n218_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n203_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G120gat), .B(G148gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(G176gat), .B(G204gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI211_X1 g062(.A(KEYINPUT12), .B(new_n227_), .C1(new_n255_), .C2(new_n218_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n251_), .A2(new_n256_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(KEYINPUT12), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n257_), .B(new_n263_), .C1(new_n266_), .C2(new_n203_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n218_), .B1(new_n243_), .B2(new_n249_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n227_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT12), .A3(new_n250_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n256_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n203_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n257_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n262_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n267_), .A2(KEYINPUT68), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT68), .B1(new_n267_), .B2(new_n276_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT13), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT13), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT69), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n285_));
  XOR2_X1   g084(.A(G183gat), .B(G211gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT76), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G127gat), .B(G155gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT74), .A3(KEYINPUT17), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(new_n269_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n290_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n289_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n302_), .B1(new_n292_), .B2(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n304_), .A2(new_n309_), .A3(KEYINPUT77), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n292_), .A2(new_n308_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n302_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n314_), .B2(new_n303_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n285_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n311_), .A3(new_n303_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n304_), .B2(new_n309_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(KEYINPUT78), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G29gat), .B(G36gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G43gat), .B(G50gat), .Z(new_n325_));
  OR3_X1    g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT15), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT15), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n218_), .B2(new_n255_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n255_), .A2(new_n218_), .A3(new_n328_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT71), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n268_), .A2(new_n331_), .A3(new_n330_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT35), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n334_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT71), .B(new_n344_), .C1(new_n333_), .C2(new_n335_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G190gat), .B(G218gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT72), .ZN(new_n348_));
  XOR2_X1   g147(.A(G134gat), .B(G162gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(KEYINPUT36), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n343_), .A2(new_n351_), .A3(new_n345_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n353_), .A2(new_n354_), .B1(KEYINPUT36), .B2(new_n350_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT37), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n350_), .A2(KEYINPUT36), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n343_), .A2(new_n351_), .A3(new_n345_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n351_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT37), .B1(new_n361_), .B2(KEYINPUT73), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n320_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT79), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  INV_X1    g167(.A(G43gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(G169gat), .B2(G176gat), .ZN(new_n376_));
  NOR3_X1   g175(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT26), .B(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT81), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n378_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n372_), .B(KEYINPUT23), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(G183gat), .B2(G190gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G169gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT82), .B(G15gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n394_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n371_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n371_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G134gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G127gat), .ZN(new_n405_));
  INV_X1    g204(.A(G127gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G134gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n407_), .A3(KEYINPUT83), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT83), .B1(new_n405_), .B2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n403_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n406_), .A2(G134gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n404_), .A2(G127gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n408_), .A3(new_n402_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT31), .ZN(new_n418_));
  OR4_X1    g217(.A1(KEYINPUT84), .A2(new_n398_), .A3(new_n401_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n401_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n400_), .B1(new_n399_), .B2(new_n395_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT84), .B1(new_n398_), .B2(new_n401_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n418_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n419_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428_));
  INV_X1    g227(.A(G141gat), .ZN(new_n429_));
  INV_X1    g228(.A(G148gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .A4(KEYINPUT85), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n432_));
  OAI22_X1  g231(.A1(new_n432_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G141gat), .A2(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT2), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n431_), .A2(new_n433_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n429_), .A2(new_n430_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n434_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT1), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n439_), .A2(new_n446_), .A3(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n427_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(G197gat), .A2(G204gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G197gat), .A2(G204gat), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G211gat), .B(G218gat), .Z(new_n454_));
  NAND4_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT87), .A4(KEYINPUT21), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(KEYINPUT21), .A3(new_n452_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G211gat), .B(G218gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n457_), .A2(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n451_), .A2(new_n452_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT21), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G228gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT86), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n450_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT88), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n459_), .A2(new_n455_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n473_));
  OAI211_X1 g272(.A(G228gat), .B(G233gat), .C1(new_n473_), .C2(new_n449_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n450_), .A2(new_n466_), .A3(new_n475_), .A4(new_n468_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n438_), .A2(new_n441_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n427_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G22gat), .B(G50gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT28), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n481_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(new_n474_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n473_), .A2(new_n449_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n475_), .B1(new_n486_), .B2(new_n468_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n471_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n479_), .A2(new_n484_), .B1(new_n477_), .B2(new_n488_), .ZN(new_n489_));
  AND4_X1   g288(.A1(KEYINPUT89), .A2(new_n488_), .A3(new_n477_), .A4(new_n484_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G85gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT0), .B(G57gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT4), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n442_), .A2(new_n448_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n416_), .A3(new_n411_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n409_), .A2(new_n403_), .A3(new_n410_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n402_), .B1(new_n415_), .B2(new_n408_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n480_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n498_), .A2(KEYINPUT93), .A3(new_n416_), .A4(new_n411_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n497_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n499_), .B2(KEYINPUT4), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n496_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT98), .ZN(new_n513_));
  INV_X1    g312(.A(new_n511_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(new_n495_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n375_), .ZN(new_n517_));
  INV_X1    g316(.A(G169gat), .ZN(new_n518_));
  INV_X1    g317(.A(G176gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n377_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n386_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n380_), .B(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n524_), .B2(new_n379_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n387_), .A2(new_n389_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n466_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n473_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(KEYINPUT20), .ZN(new_n529_));
  NAND3_X1  g328(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT90), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n391_), .A2(new_n466_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n533_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT20), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT26), .B(G190gat), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n523_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n380_), .A2(KEYINPUT91), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n379_), .A3(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n541_), .A2(new_n378_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n537_), .B1(new_n542_), .B2(new_n473_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n529_), .A2(new_n534_), .B1(new_n535_), .B2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G8gat), .B(G36gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G64gat), .B(G92gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT32), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n542_), .B2(new_n473_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n535_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n533_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n541_), .A2(new_n378_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n390_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n559_), .B2(new_n466_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n534_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n528_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n550_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n551_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n544_), .A2(KEYINPUT96), .A3(new_n550_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT98), .B(new_n496_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n516_), .A2(new_n565_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT94), .B1(KEYINPUT95), .B2(KEYINPUT33), .ZN(new_n569_));
  NOR2_X1   g368(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n515_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n549_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n561_), .B1(new_n560_), .B2(new_n528_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n543_), .A2(new_n535_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n529_), .A2(new_n534_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n543_), .A2(new_n535_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n549_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n504_), .A2(new_n505_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT4), .ZN(new_n581_));
  INV_X1    g380(.A(new_n509_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n511_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n570_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n569_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n583_), .A2(new_n495_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n495_), .B1(new_n580_), .B2(new_n508_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n507_), .B1(new_n499_), .B2(KEYINPUT4), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n506_), .B2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n571_), .A2(new_n579_), .A3(new_n586_), .A4(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n491_), .B1(new_n568_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n516_), .A2(new_n567_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n575_), .A2(new_n578_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT27), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n562_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n536_), .B1(new_n554_), .B2(new_n535_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n572_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n593_), .A2(new_n594_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n592_), .A2(new_n491_), .A3(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n426_), .B1(new_n591_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT99), .ZN(new_n602_));
  INV_X1    g401(.A(new_n592_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n426_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n491_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n599_), .A2(KEYINPUT100), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n599_), .A2(KEYINPUT100), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n604_), .B(new_n605_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n426_), .C1(new_n591_), .C2(new_n600_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n332_), .A2(new_n299_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n299_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n328_), .A2(new_n299_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n615_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n616_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n613_), .A2(new_n618_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT80), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n624_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n612_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n284_), .A2(new_n367_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n294_), .A3(new_n603_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT101), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT101), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n635_), .A2(KEYINPUT38), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT38), .B1(new_n635_), .B2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n611_), .A2(new_n355_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n310_), .A2(new_n315_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n283_), .A2(new_n641_), .A3(new_n629_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT102), .B1(new_n639_), .B2(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n294_), .B1(new_n647_), .B2(new_n603_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n637_), .A2(new_n638_), .A3(new_n648_), .ZN(G1324gat));
  OR2_X1    g448(.A1(new_n607_), .A2(new_n606_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n633_), .A2(new_n295_), .A3(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT39), .B(new_n295_), .C1(new_n643_), .C2(new_n651_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n643_), .A2(new_n651_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g457(.A(new_n647_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n426_), .ZN(new_n660_));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n660_), .A2(KEYINPUT103), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT103), .B1(new_n660_), .B2(new_n661_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n426_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n633_), .A2(new_n661_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n662_), .A2(KEYINPUT41), .A3(new_n663_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n666_), .A2(new_n668_), .A3(new_n669_), .ZN(G1326gat));
  OR3_X1    g469(.A1(new_n632_), .A2(G22gat), .A3(new_n605_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G22gat), .B1(new_n659_), .B2(new_n605_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT42), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(KEYINPUT42), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1327gat));
  AND3_X1   g474(.A1(new_n317_), .A2(new_n318_), .A3(KEYINPUT78), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT78), .B1(new_n317_), .B2(new_n318_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT104), .B1(new_n678_), .B2(new_n355_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n320_), .A2(new_n680_), .A3(new_n363_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n679_), .A2(new_n681_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n631_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n603_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n283_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(new_n678_), .A3(new_n630_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n363_), .B(new_n358_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n601_), .A2(KEYINPUT99), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n610_), .A2(new_n608_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n688_), .B(new_n689_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n688_), .B1(new_n611_), .B2(new_n689_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n687_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n687_), .B(KEYINPUT44), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n603_), .A2(G29gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n685_), .B1(new_n699_), .B2(new_n700_), .ZN(G1328gat));
  NOR2_X1   g500(.A1(new_n650_), .A2(G36gat), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n682_), .A2(new_n611_), .A3(new_n629_), .A4(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n697_), .A2(new_n651_), .A3(new_n698_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(G36gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT46), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT107), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n705_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT46), .B1(new_n713_), .B2(KEYINPUT105), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT105), .B(new_n705_), .C1(new_n706_), .C2(G36gat), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n710_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n707_), .B2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(KEYINPUT106), .A3(new_n715_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n709_), .B1(new_n717_), .B2(new_n721_), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n699_), .A2(G43gat), .A3(new_n667_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n369_), .B1(new_n683_), .B2(new_n426_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n684_), .B2(new_n491_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n491_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n699_), .B2(new_n728_), .ZN(G1331gat));
  NOR4_X1   g528(.A1(new_n284_), .A2(new_n320_), .A3(new_n629_), .A4(new_n639_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT111), .B(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n603_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n611_), .A2(new_n630_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT109), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n367_), .A2(new_n686_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT108), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT108), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n603_), .B(new_n734_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(KEYINPUT110), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT110), .B1(new_n738_), .B2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n732_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT112), .B(new_n732_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n730_), .A2(new_n651_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G64gat), .ZN(new_n749_));
  INV_X1    g548(.A(G64gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT48), .B(new_n750_), .C1(new_n730_), .C2(new_n651_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n651_), .A2(new_n750_), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n749_), .A2(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT113), .Z(G1333gat));
  INV_X1    g554(.A(new_n730_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G71gat), .B1(new_n756_), .B2(new_n426_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n426_), .A2(G71gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n752_), .B2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n756_), .B2(new_n605_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT50), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n605_), .A2(G78gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n752_), .B2(new_n763_), .ZN(G1335gat));
  OR2_X1    g563(.A1(new_n693_), .A2(new_n694_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n283_), .A2(new_n678_), .A3(new_n629_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n592_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n284_), .B1(new_n681_), .B2(new_n679_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n734_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n603_), .A2(new_n209_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1336gat));
  OAI21_X1  g571(.A(G92gat), .B1(new_n767_), .B2(new_n650_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n651_), .A2(new_n210_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n770_), .B2(new_n774_), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n767_), .B2(new_n426_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n667_), .A2(new_n213_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n770_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n491_), .A3(new_n766_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n491_), .A2(new_n214_), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n782_), .A2(new_n783_), .B1(new_n770_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n650_), .A2(new_n605_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n667_), .A2(new_n603_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n629_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n366_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(new_n366_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n271_), .A2(new_n273_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n202_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n271_), .A2(new_n203_), .A3(new_n273_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(KEYINPUT55), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n801_), .A3(new_n202_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n262_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n263_), .A2(new_n804_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(new_n802_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n800_), .A2(KEYINPUT114), .A3(new_n802_), .A4(new_n806_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n805_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n629_), .A2(new_n267_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n622_), .A2(new_n628_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n613_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n620_), .A2(new_n616_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n627_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n277_), .A2(new_n278_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n813_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n355_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n267_), .B1(new_n817_), .B2(new_n814_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n365_), .B(new_n359_), .C1(new_n824_), .C2(KEYINPUT58), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(new_n823_), .C1(new_n805_), .C2(new_n807_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n819_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n355_), .A2(KEYINPUT57), .ZN(new_n829_));
  OAI22_X1  g628(.A1(new_n825_), .A2(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n320_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n796_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n824_), .A2(KEYINPUT58), .ZN(new_n834_));
  INV_X1    g633(.A(new_n827_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n689_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n828_), .B2(new_n363_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n829_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n821_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT117), .A3(new_n320_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n791_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n836_), .A2(new_n838_), .A3(new_n840_), .A4(KEYINPUT115), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n640_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n796_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n789_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n843_), .B1(new_n850_), .B2(KEYINPUT59), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n630_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n630_), .A2(G113gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n850_), .B2(new_n854_), .ZN(G1340gat));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n284_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n851_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n850_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n283_), .B2(KEYINPUT60), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n857_), .B2(KEYINPUT60), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n856_), .B1(new_n859_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n641_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n796_), .B1(new_n869_), .B2(new_n846_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n789_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT59), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n843_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n858_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G120gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT119), .A3(new_n866_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n868_), .A2(new_n876_), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n852_), .B2(new_n640_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n860_), .A2(new_n406_), .A3(new_n678_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1342gat));
  INV_X1    g679(.A(new_n689_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G134gat), .B1(new_n852_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n860_), .A2(new_n404_), .A3(new_n363_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1343gat));
  NOR4_X1   g683(.A1(new_n651_), .A2(new_n667_), .A3(new_n605_), .A4(new_n592_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n849_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n629_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n849_), .A2(new_n885_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT121), .B1(new_n889_), .B2(new_n630_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT120), .B(G141gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n891_), .B(new_n893_), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n889_), .A2(new_n284_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n430_), .ZN(G1345gat));
  NAND3_X1  g695(.A1(new_n886_), .A2(KEYINPUT122), .A3(new_n678_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n889_), .B2(new_n320_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n889_), .B2(new_n355_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT123), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n889_), .A2(new_n903_), .A3(new_n881_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1347gat));
  NAND2_X1  g706(.A1(new_n833_), .A2(new_n842_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n650_), .A2(new_n426_), .A3(new_n603_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n909_), .A2(new_n605_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT124), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n910_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT22), .B(G169gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n629_), .A3(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n518_), .B1(new_n911_), .B2(new_n629_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n920_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n918_), .B1(new_n921_), .B2(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n870_), .A2(new_n491_), .ZN(new_n924_));
  AND4_X1   g723(.A1(G176gat), .A2(new_n924_), .A3(new_n858_), .A4(new_n909_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n916_), .A2(new_n686_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n519_), .ZN(G1349gat));
  AND2_X1   g726(.A1(new_n909_), .A2(new_n678_), .ZN(new_n928_));
  AOI21_X1  g727(.A(G183gat), .B1(new_n924_), .B2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n640_), .A2(new_n379_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n916_), .B2(new_n930_), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n916_), .A2(new_n363_), .A3(new_n524_), .ZN(new_n932_));
  INV_X1    g731(.A(G190gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n881_), .B1(new_n912_), .B2(new_n915_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1351gat));
  NAND3_X1  g734(.A1(new_n426_), .A2(new_n491_), .A3(new_n592_), .ZN(new_n936_));
  XOR2_X1   g735(.A(new_n936_), .B(KEYINPUT125), .Z(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n650_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n849_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT126), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n849_), .A2(new_n941_), .A3(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(KEYINPUT127), .B(G197gat), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n943_), .A2(new_n629_), .A3(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n943_), .B2(new_n629_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1352gat));
  INV_X1    g746(.A(new_n943_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G204gat), .B1(new_n948_), .B2(new_n284_), .ZN(new_n949_));
  INV_X1    g748(.A(G204gat), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n943_), .A2(new_n950_), .A3(new_n858_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n951_), .ZN(G1353gat));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n640_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n943_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n943_), .B2(new_n955_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n948_), .B2(new_n881_), .ZN(new_n959_));
  INV_X1    g758(.A(G218gat), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n943_), .A2(new_n960_), .A3(new_n363_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1355gat));
endmodule


