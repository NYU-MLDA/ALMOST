//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT38), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G71gat), .B(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G227gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(G15gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G43gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n208_), .B(G15gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(G43gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT30), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(G43gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n211_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(new_n206_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n215_), .B2(new_n219_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  INV_X1    g025(.A(G176gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT83), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(KEYINPUT83), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT84), .B1(new_n232_), .B2(KEYINPUT23), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(KEYINPUT23), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(KEYINPUT84), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n229_), .B(new_n230_), .C1(new_n231_), .C2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT25), .B(G183gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT26), .B(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G169gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n227_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT24), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n239_), .A2(new_n234_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT85), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n223_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n223_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT31), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT31), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n248_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n223_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n256_), .B2(new_n249_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G127gat), .B(G134gat), .Z(new_n258_));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n252_), .A2(new_n257_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT31), .B1(new_n250_), .B2(new_n251_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(new_n253_), .A3(new_n249_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n205_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G197gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n267_), .A2(G204gat), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT21), .ZN(new_n272_));
  XOR2_X1   g071(.A(G211gat), .B(G218gat), .Z(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n270_), .B(KEYINPUT89), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n268_), .B(KEYINPUT90), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT21), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n273_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  OR3_X1    g084(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n282_), .A2(KEYINPUT1), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n297_), .A3(new_n281_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G141gat), .B(G148gat), .Z(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT87), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT87), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n294_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n280_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(G228gat), .A2(G233gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n280_), .B(new_n309_), .C1(new_n303_), .C2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT92), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G22gat), .B(G50gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT28), .B1(new_n302_), .B2(KEYINPUT29), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n301_), .A2(new_n300_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n310_), .A4(new_n294_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n315_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(new_n319_), .A3(new_n315_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n313_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n324_), .A2(new_n312_), .A3(new_n320_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n308_), .B(new_n311_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(KEYINPUT92), .B(new_n312_), .C1(new_n324_), .C2(new_n320_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n308_), .A2(new_n311_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n322_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n327_), .B(new_n328_), .C1(new_n312_), .C2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n261_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n263_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT86), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n266_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n326_), .A2(new_n330_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n234_), .B1(G183gat), .B2(G190gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n228_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n239_), .A2(new_n243_), .A3(new_n242_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n235_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT94), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(KEYINPUT94), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n341_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n339_), .B1(new_n347_), .B2(new_n280_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n280_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n246_), .A2(new_n349_), .A3(new_n248_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n235_), .A2(new_n342_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n358_), .A2(new_n344_), .B1(new_n228_), .B2(new_n340_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n339_), .B(new_n354_), .C1(new_n359_), .C2(new_n349_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n349_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND3_X1  g166(.A1(new_n355_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n354_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT20), .B(new_n370_), .C1(new_n347_), .C2(new_n280_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(new_n361_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n369_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n341_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n280_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n354_), .B1(new_n361_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n369_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT27), .A3(new_n368_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n302_), .A2(new_n260_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n261_), .A2(new_n317_), .A3(new_n294_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT95), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n303_), .A2(KEYINPUT95), .A3(new_n261_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n385_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G57gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n388_), .A2(new_n391_), .A3(new_n389_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n395_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n395_), .B2(new_n401_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n384_), .A2(new_n405_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n262_), .A2(new_n265_), .A3(new_n205_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT86), .B1(new_n332_), .B2(new_n333_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n331_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n371_), .A2(new_n373_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n411_));
  MUX2_X1   g210(.A(new_n381_), .B(new_n410_), .S(new_n411_), .Z(new_n412_));
  AND3_X1   g211(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n388_), .A2(new_n392_), .A3(new_n389_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT33), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n400_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n395_), .A2(new_n417_), .A3(new_n401_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n416_), .A2(new_n368_), .A3(new_n374_), .A4(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n403_), .A2(KEYINPUT33), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n412_), .A2(new_n404_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n338_), .A2(new_n406_), .B1(new_n409_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n423_));
  XOR2_X1   g222(.A(G29gat), .B(G36gat), .Z(new_n424_));
  XOR2_X1   g223(.A(G43gat), .B(G50gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT15), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G22gat), .ZN(new_n428_));
  INV_X1    g227(.A(G1gat), .ZN(new_n429_));
  INV_X1    g228(.A(G8gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT14), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G8gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n426_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n436_), .A2(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G229gat), .A2(G233gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n436_), .B(new_n434_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n438_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G113gat), .B(G141gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G169gat), .B(G197gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n443_), .A2(new_n447_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n423_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(KEYINPUT82), .A3(new_n448_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n422_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G190gat), .B(G218gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT78), .ZN(new_n457_));
  XOR2_X1   g256(.A(G134gat), .B(G162gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n463_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT64), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n467_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT9), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT64), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  AND3_X1   g277(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT10), .B(G99gat), .Z(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  AOI211_X1 g280(.A(new_n478_), .B(new_n479_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n479_), .A2(new_n478_), .ZN(new_n484_));
  OR3_X1    g283(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT65), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT66), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n483_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n462_), .B1(new_n496_), .B2(new_n436_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n478_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n485_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n488_), .A2(new_n489_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n492_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT8), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n503_), .A2(new_n493_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT76), .A3(new_n426_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(KEYINPUT72), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT72), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n483_), .B(new_n508_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n427_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n506_), .A2(new_n510_), .A3(KEYINPUT77), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT35), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n506_), .A2(new_n511_), .A3(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n512_), .A2(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n512_), .A2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n459_), .A2(new_n460_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n461_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT37), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n525_), .B2(KEYINPUT80), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n523_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n532_));
  OAI22_X1  g331(.A1(new_n531_), .A2(new_n532_), .B1(new_n460_), .B2(new_n459_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT80), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT37), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539_));
  AND2_X1   g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n434_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(G57gat), .ZN(new_n544_));
  INV_X1    g343(.A(G57gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G64gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n546_), .A3(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT68), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n544_), .A2(new_n546_), .A3(new_n549_), .A4(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n544_), .A2(new_n546_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT11), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G78gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT11), .B1(new_n544_), .B2(new_n546_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT67), .B1(new_n559_), .B2(new_n556_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n549_), .B1(new_n562_), .B2(KEYINPUT11), .ZN(new_n563_));
  INV_X1    g362(.A(new_n550_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n555_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n559_), .A2(KEYINPUT67), .A3(new_n556_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n542_), .B1(new_n561_), .B2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT16), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n551_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n551_), .B1(new_n560_), .B2(new_n558_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n541_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  OR4_X1    g375(.A1(new_n539_), .A2(new_n569_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n573_), .B(KEYINPUT17), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n568_), .A2(KEYINPUT69), .A3(new_n561_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n542_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n541_), .A2(new_n581_), .A3(new_n580_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n578_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT81), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n586_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n577_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n538_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n455_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n580_), .A2(new_n581_), .A3(new_n504_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n568_), .A2(KEYINPUT69), .A3(new_n561_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT69), .B1(new_n568_), .B2(new_n561_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n496_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT70), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n504_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n594_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n592_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n600_), .B1(new_n582_), .B2(new_n496_), .ZN(new_n605_));
  AOI211_X1 g404(.A(KEYINPUT70), .B(new_n504_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n593_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n603_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(KEYINPUT71), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n568_), .B2(new_n561_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n507_), .A2(new_n509_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n599_), .B2(KEYINPUT12), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n593_), .A2(new_n603_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n593_), .A2(KEYINPUT73), .A3(new_n603_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n610_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT5), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n610_), .A2(new_n620_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(KEYINPUT13), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n610_), .B2(new_n620_), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n619_), .B(new_n625_), .C1(new_n604_), .C2(new_n609_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT74), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n591_), .A2(new_n429_), .A3(new_n405_), .A4(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n202_), .A2(new_n203_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n204_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n589_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n454_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n643_), .A2(KEYINPUT96), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n533_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n422_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(KEYINPUT96), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n644_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n404_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n640_), .B(new_n652_), .C1(new_n204_), .C2(new_n638_), .ZN(G1324gat));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT101), .Z(new_n655_));
  NAND4_X1  g454(.A1(new_n644_), .A2(new_n384_), .A3(new_n648_), .A4(new_n649_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(G8gat), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n656_), .B2(G8gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT39), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n658_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n636_), .A2(new_n591_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n384_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n666_), .A2(G8gat), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n655_), .B1(new_n665_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n655_), .ZN(new_n671_));
  AOI211_X1 g470(.A(new_n668_), .B(new_n671_), .C1(new_n661_), .C2(new_n664_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1325gat));
  NOR2_X1   g472(.A1(new_n407_), .A2(new_n408_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n209_), .B1(new_n650_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT41), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n209_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n666_), .B2(new_n678_), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n650_), .A2(new_n331_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G22gat), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT103), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT103), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n336_), .A2(G22gat), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT104), .Z(new_n688_));
  OAI22_X1  g487(.A1(new_n685_), .A2(new_n686_), .B1(new_n666_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n634_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n641_), .A3(new_n454_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n338_), .A2(new_n406_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n409_), .A2(new_n421_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(KEYINPUT105), .A3(new_n695_), .A4(new_n538_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n422_), .B2(new_n537_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n422_), .A2(new_n537_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n699_), .B2(new_n695_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n691_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n694_), .A2(new_n538_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n697_), .A3(new_n696_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n708_), .A3(new_n405_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G29gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n527_), .A2(new_n641_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n455_), .A2(new_n634_), .A3(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n404_), .A2(G29gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT106), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n703_), .A2(new_n708_), .A3(new_n384_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  INV_X1    g518(.A(G36gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n720_), .A3(new_n384_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT45), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT107), .B(new_n717_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n717_), .A2(KEYINPUT107), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n717_), .A2(KEYINPUT107), .ZN(new_n725_));
  AND4_X1   g524(.A1(new_n724_), .A2(new_n719_), .A3(new_n725_), .A4(new_n722_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1329gat));
  NOR2_X1   g526(.A1(new_n262_), .A2(new_n265_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n211_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n703_), .A2(new_n708_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT108), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n703_), .A2(new_n708_), .A3(new_n732_), .A4(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n712_), .A2(new_n675_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n211_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n731_), .A2(new_n738_), .A3(new_n733_), .A4(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1330gat));
  INV_X1    g539(.A(G50gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n703_), .A2(new_n708_), .A3(new_n331_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(KEYINPUT109), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(KEYINPUT109), .B2(new_n742_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n712_), .A2(new_n741_), .A3(new_n331_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n642_), .A2(new_n589_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n635_), .A2(new_n648_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n404_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n422_), .A2(new_n642_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(new_n690_), .A3(new_n590_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n545_), .A3(new_n405_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1332gat));
  NAND3_X1  g552(.A1(new_n751_), .A2(new_n543_), .A3(new_n384_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G64gat), .B1(new_n748_), .B2(new_n667_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT111), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT111), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n758_));
  AND3_X1   g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n754_), .B1(new_n759_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n748_), .B2(new_n674_), .ZN(new_n762_));
  XOR2_X1   g561(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n751_), .A2(new_n765_), .A3(new_n675_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1334gat));
  OAI21_X1  g566(.A(G78gat), .B1(new_n748_), .B2(new_n336_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT50), .ZN(new_n769_));
  INV_X1    g568(.A(G78gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n751_), .A2(new_n770_), .A3(new_n331_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n634_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n707_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n404_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n635_), .A2(new_n750_), .A3(new_n711_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n464_), .A3(new_n405_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1336gat));
  OAI21_X1  g577(.A(G92gat), .B1(new_n774_), .B2(new_n667_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n465_), .A3(new_n384_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n774_), .B2(new_n674_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n776_), .B(new_n480_), .C1(new_n262_), .C2(new_n265_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(KEYINPUT113), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n784_), .B(new_n786_), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n776_), .A2(new_n481_), .A3(new_n331_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n331_), .B(new_n773_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n707_), .A2(KEYINPUT114), .A3(new_n331_), .A4(new_n773_), .ZN(new_n793_));
  AND4_X1   g592(.A1(new_n789_), .A2(new_n792_), .A3(new_n793_), .A4(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n481_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n789_), .B1(new_n795_), .B2(new_n793_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n788_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n788_), .C1(new_n794_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NAND3_X1  g600(.A1(new_n435_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n446_), .B1(new_n440_), .B2(new_n438_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n450_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT119), .B(new_n804_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n632_), .A2(new_n454_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n593_), .A2(KEYINPUT73), .A3(new_n603_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT73), .B1(new_n593_), .B2(new_n603_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n814_), .B2(new_n614_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n614_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(KEYINPUT55), .C1(new_n813_), .C2(new_n812_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n613_), .B(new_n593_), .C1(new_n599_), .C2(KEYINPUT12), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n608_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n821_), .A3(new_n608_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n815_), .A2(new_n817_), .A3(new_n820_), .A4(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n625_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n823_), .B2(new_n625_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n810_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n810_), .B(new_n829_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n809_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n533_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n804_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT120), .B1(new_n632_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n628_), .A2(new_n837_), .A3(new_n804_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n625_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n836_), .B(new_n838_), .C1(new_n824_), .C2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n537_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n824_), .A2(new_n839_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(KEYINPUT58), .A3(new_n838_), .A4(new_n836_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n834_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n831_), .B2(new_n527_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n589_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n629_), .A2(new_n633_), .A3(new_n747_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT115), .B1(new_n538_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n634_), .A2(new_n851_), .A3(new_n537_), .A4(new_n747_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n852_), .A3(KEYINPUT54), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT115), .B(new_n854_), .C1(new_n538_), .C2(new_n849_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n384_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n337_), .A2(new_n404_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT59), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n831_), .A2(new_n527_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n832_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n831_), .A2(new_n833_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n641_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n667_), .B(new_n859_), .C1(new_n864_), .C2(new_n856_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n860_), .A2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n454_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n865_), .A2(G113gat), .A3(new_n454_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1340gat));
  OAI21_X1  g670(.A(G120gat), .B1(new_n868_), .B2(new_n636_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n865_), .ZN(new_n873_));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n634_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n873_), .B(new_n875_), .C1(KEYINPUT60), .C2(new_n874_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n876_), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n868_), .B2(new_n589_), .ZN(new_n878_));
  OR3_X1    g677(.A1(new_n865_), .A2(G127gat), .A3(new_n589_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n537_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n865_), .B2(new_n646_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(KEYINPUT121), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886_));
  INV_X1    g685(.A(new_n882_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n858_), .A2(KEYINPUT59), .A3(new_n859_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n865_), .A2(new_n866_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n884_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n886_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n885_), .A2(new_n892_), .ZN(G1343gat));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n335_), .A2(new_n404_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n858_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n667_), .B(new_n895_), .C1(new_n864_), .C2(new_n856_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT122), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n454_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n288_), .ZN(G1344gat));
  AOI21_X1  g699(.A(new_n636_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n289_), .ZN(G1345gat));
  AOI21_X1  g701(.A(new_n589_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT123), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n903_), .B(new_n906_), .ZN(G1346gat));
  NAND2_X1  g706(.A1(new_n896_), .A2(new_n898_), .ZN(new_n908_));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(new_n647_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n537_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(new_n911_), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n848_), .A2(new_n857_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n384_), .A2(new_n404_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n914_), .A2(new_n674_), .A3(new_n331_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916_), .B2(new_n454_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n916_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n642_), .A3(new_n226_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n918_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n916_), .B2(new_n636_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n690_), .A2(new_n227_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n916_), .B2(new_n925_), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n916_), .A2(new_n589_), .ZN(new_n927_));
  MUX2_X1   g726(.A(G183gat), .B(new_n237_), .S(new_n927_), .Z(G1350gat));
  NAND4_X1  g727(.A1(new_n913_), .A2(new_n238_), .A3(new_n647_), .A4(new_n915_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n538_), .B(new_n915_), .C1(new_n864_), .C2(new_n856_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n930_), .A2(new_n931_), .A3(G190gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(G190gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n929_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT125), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n936_), .B(new_n929_), .C1(new_n932_), .C2(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n864_), .A2(new_n856_), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n914_), .A2(new_n335_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n642_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n635_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G204gat), .ZN(G1353gat));
  OR3_X1    g744(.A1(new_n939_), .A2(new_n589_), .A3(new_n940_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n946_), .A2(KEYINPUT127), .A3(new_n947_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT63), .B(G211gat), .Z(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n952_), .B1(new_n946_), .B2(new_n954_), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n941_), .A2(KEYINPUT126), .A3(new_n641_), .A4(new_n953_), .ZN(new_n956_));
  AOI22_X1  g755(.A1(new_n950_), .A2(new_n951_), .B1(new_n955_), .B2(new_n956_), .ZN(G1354gat));
  INV_X1    g756(.A(G218gat), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n941_), .A2(new_n958_), .A3(new_n647_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n939_), .A2(new_n537_), .A3(new_n940_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n958_), .B2(new_n960_), .ZN(G1355gat));
endmodule


