//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT94), .B(G197gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(G204gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(G197gat), .B2(G204gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n209_), .A2(new_n213_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n208_), .A2(new_n215_), .B1(new_n206_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT1), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT92), .Z(new_n223_));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(KEYINPUT1), .B2(new_n221_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n218_), .B(new_n220_), .C1(new_n223_), .C2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n219_), .B(KEYINPUT3), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n218_), .B(KEYINPUT2), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT93), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(new_n221_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n217_), .B1(new_n233_), .B2(KEYINPUT29), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT95), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(G228gat), .B2(G233gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(G78gat), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n234_), .A2(G78gat), .A3(new_n236_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n203_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n238_), .A2(new_n203_), .A3(new_n239_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n202_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT28), .Z(new_n249_));
  NAND3_X1  g048(.A1(new_n235_), .A2(G228gat), .A3(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G64gat), .B(G92gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT99), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT19), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G169gat), .B(G176gat), .ZN(new_n271_));
  INV_X1    g070(.A(G183gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT25), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276_));
  AOI22_X1  g075(.A1(KEYINPUT83), .A2(new_n273_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(KEYINPUT83), .B2(new_n273_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n272_), .A2(KEYINPUT25), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n279_), .B(new_n280_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n281_));
  OAI221_X1 g080(.A(new_n270_), .B1(new_n268_), .B2(new_n271_), .C1(new_n278_), .C2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n265_), .B2(KEYINPUT23), .ZN(new_n286_));
  INV_X1    g085(.A(new_n267_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n284_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT86), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n217_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT96), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT20), .ZN(new_n295_));
  INV_X1    g094(.A(new_n217_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n271_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n269_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n279_), .A2(new_n273_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n280_), .A2(new_n275_), .ZN(new_n302_));
  OAI221_X1 g101(.A(new_n299_), .B1(new_n300_), .B2(new_n298_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n267_), .A2(new_n289_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n304_), .A2(KEYINPUT98), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n284_), .B1(new_n304_), .B2(KEYINPUT98), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n303_), .A2(new_n288_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n296_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n295_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n294_), .B1(new_n293_), .B2(KEYINPUT20), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n262_), .B(new_n264_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n296_), .A2(new_n307_), .ZN(new_n312_));
  OAI211_X1 g111(.A(KEYINPUT20), .B(new_n312_), .C1(new_n292_), .C2(new_n217_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n313_), .A2(new_n264_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n293_), .A2(KEYINPUT20), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT96), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n308_), .A3(new_n295_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n262_), .B1(new_n318_), .B2(new_n264_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n261_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n264_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT99), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n322_), .A2(new_n260_), .A3(new_n314_), .A4(new_n311_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT27), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT27), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n313_), .A2(new_n264_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n318_), .B2(new_n264_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n327_), .B2(new_n261_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n328_), .A2(new_n323_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n233_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n233_), .A2(new_n335_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(KEYINPUT4), .C1(KEYINPUT100), .C2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT100), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n233_), .A2(new_n339_), .A3(new_n340_), .A4(new_n335_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n330_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G85gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT0), .B(G57gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  AOI22_X1  g145(.A1(new_n336_), .A2(new_n337_), .B1(G225gat), .B2(G233gat), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n342_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT87), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT30), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT31), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n335_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT88), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G99gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(G71gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G99gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(KEYINPUT88), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n354_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n354_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n292_), .B(KEYINPUT91), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n351_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NOR4_X1   g173(.A1(new_n256_), .A2(new_n324_), .A3(new_n329_), .A4(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n327_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n322_), .A2(new_n314_), .A3(new_n311_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n350_), .B(new_n377_), .C1(new_n378_), .C2(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n320_), .A2(new_n323_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n338_), .A2(new_n330_), .A3(new_n341_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n346_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT101), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n336_), .A2(new_n384_), .A3(new_n337_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n330_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT33), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  MUX2_X1   g187(.A(KEYINPUT33), .B(new_n388_), .S(new_n349_), .Z(new_n389_));
  OAI21_X1  g188(.A(new_n379_), .B1(new_n380_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n255_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n255_), .A2(new_n350_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n380_), .A2(new_n325_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n328_), .A2(new_n323_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n372_), .A2(new_n373_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n375_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G29gat), .B(G36gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G43gat), .B(G50gat), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n400_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G15gat), .ZN(new_n404_));
  INV_X1    g203(.A(G22gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G15gat), .A2(G22gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G1gat), .A2(G8gat), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n406_), .A2(new_n407_), .B1(KEYINPUT14), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(G15gat), .A2(G22gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G15gat), .A2(G22gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n408_), .A2(KEYINPUT14), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT78), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n411_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n411_), .B2(new_n416_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G1gat), .B(G8gat), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n411_), .A2(new_n416_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT79), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n411_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n403_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n403_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G229gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n401_), .A2(KEYINPUT15), .A3(new_n402_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT15), .B1(new_n401_), .B2(new_n402_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n428_), .A2(new_n429_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n427_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G113gat), .B(G141gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT82), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G169gat), .B(G197gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n435_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n422_), .A2(new_n426_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G231gat), .A2(G233gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT80), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n450_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT70), .B(G71gat), .ZN(new_n454_));
  INV_X1    g253(.A(G78gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G57gat), .B(G64gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT11), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n454_), .A2(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n455_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n458_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n457_), .A2(KEYINPUT11), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n460_), .B(new_n461_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n453_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G127gat), .B(G155gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT16), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G183gat), .B(G211gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT17), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n468_), .A2(new_n475_), .A3(new_n472_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(new_n477_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n474_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT34), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT35), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT64), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT64), .B1(new_n488_), .B2(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n203_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT66), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT65), .B(G92gat), .ZN(new_n495_));
  INV_X1    g294(.A(G85gat), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT9), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n493_), .A2(new_n494_), .A3(new_n498_), .A4(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT10), .B(G99gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(G106gat), .B1(new_n512_), .B2(new_n490_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n503_), .B(new_n507_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT66), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT67), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n505_), .A2(new_n525_), .A3(new_n506_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(KEYINPUT68), .A3(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n517_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n503_), .A2(KEYINPUT69), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n500_), .A2(new_n502_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n505_), .A2(new_n506_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n525_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n516_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n540_), .A2(new_n438_), .B1(new_n485_), .B2(new_n484_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT68), .B1(new_n524_), .B2(new_n527_), .ZN(new_n543_));
  AOI211_X1 g342(.A(new_n529_), .B(new_n526_), .C1(new_n518_), .C2(new_n523_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n538_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT8), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n545_), .A2(new_n547_), .B1(new_n515_), .B2(new_n509_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n403_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n542_), .B1(new_n541_), .B2(new_n549_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n487_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n540_), .A2(new_n438_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n484_), .A2(new_n485_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT75), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(new_n486_), .A3(new_n550_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT36), .Z(new_n562_));
  NAND3_X1  g361(.A1(new_n553_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n566_), .B2(KEYINPUT76), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n551_), .A2(new_n552_), .A3(new_n487_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n486_), .B1(new_n557_), .B2(new_n550_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT76), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n562_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n481_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n564_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT77), .A3(new_n563_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT77), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n576_), .A3(new_n562_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT37), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n480_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT12), .B1(new_n548_), .B2(new_n465_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n540_), .A2(new_n582_), .A3(new_n466_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n516_), .B(new_n465_), .C1(new_n532_), .C2(new_n539_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(KEYINPUT72), .A3(new_n586_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n584_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(KEYINPUT71), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n540_), .A2(new_n466_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n545_), .A2(new_n547_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n516_), .A4(new_n465_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n586_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT74), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n591_), .A2(new_n599_), .A3(new_n606_), .A4(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n591_), .A2(new_n599_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n603_), .B(KEYINPUT73), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n608_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n580_), .A2(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n398_), .A2(new_n449_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n619_), .A2(G1gat), .A3(new_n351_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n396_), .A2(new_n397_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n375_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n575_), .A2(new_n577_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n480_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n616_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n449_), .ZN(new_n628_));
  AND4_X1   g427(.A1(new_n623_), .A2(new_n625_), .A3(new_n626_), .A4(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n350_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n620_), .A2(KEYINPUT38), .B1(new_n630_), .B2(G1gat), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632_));
  INV_X1    g431(.A(new_n620_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n620_), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1324gat));
  INV_X1    g438(.A(G8gat), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n324_), .A2(new_n329_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n618_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n629_), .A2(new_n642_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G8gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT39), .B(new_n640_), .C1(new_n629_), .C2(new_n642_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g448(.A(new_n397_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n404_), .B1(new_n629_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT41), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n618_), .A2(new_n404_), .A3(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  XOR2_X1   g453(.A(new_n255_), .B(KEYINPUT104), .Z(new_n655_));
  AOI21_X1  g454(.A(new_n405_), .B1(new_n629_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT42), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n618_), .A2(new_n405_), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1327gat));
  NOR2_X1   g458(.A1(new_n398_), .A2(new_n449_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n626_), .A2(new_n625_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n616_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n350_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n573_), .A2(new_n578_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n398_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n650_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT43), .B(new_n579_), .C1(new_n668_), .C2(new_n375_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n667_), .A2(new_n480_), .A3(new_n628_), .A4(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(KEYINPUT105), .A3(new_n671_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n350_), .A2(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n664_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n677_), .B2(new_n642_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n662_), .A2(G36gat), .A3(new_n641_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n672_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n676_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT105), .B1(new_n670_), .B2(new_n671_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G36gat), .B1(new_n689_), .B2(new_n641_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n684_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT46), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n685_), .A2(new_n692_), .ZN(G1329gat));
  INV_X1    g492(.A(G43gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n397_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n677_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n662_), .B2(new_n397_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT47), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(new_n700_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n663_), .B2(new_n655_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n256_), .A2(G50gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n677_), .B2(new_n704_), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n616_), .A2(new_n448_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR4_X1   g506(.A1(new_n398_), .A2(new_n624_), .A3(new_n480_), .A4(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n351_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n398_), .A2(new_n707_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n580_), .ZN(new_n712_));
  INV_X1    g511(.A(G57gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n350_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1332gat));
  INV_X1    g514(.A(G64gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n708_), .B2(new_n642_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT48), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n712_), .A2(new_n716_), .A3(new_n642_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1333gat));
  AOI21_X1  g519(.A(new_n360_), .B1(new_n708_), .B2(new_n650_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT49), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n712_), .A2(new_n360_), .A3(new_n650_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1334gat));
  AOI21_X1  g523(.A(new_n455_), .B1(new_n708_), .B2(new_n655_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT50), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n712_), .A2(new_n455_), .A3(new_n655_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1335gat));
  NAND2_X1  g527(.A1(new_n711_), .A2(new_n661_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n496_), .B1(new_n729_), .B2(new_n351_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT106), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n623_), .A2(new_n579_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n626_), .B1(new_n732_), .B2(new_n665_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n669_), .A3(new_n706_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(new_n496_), .A3(new_n351_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1336gat));
  OAI21_X1  g535(.A(new_n504_), .B1(new_n729_), .B2(new_n641_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT107), .Z(new_n738_));
  NOR3_X1   g537(.A1(new_n734_), .A2(new_n641_), .A3(new_n495_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1337gat));
  AOI211_X1 g539(.A(new_n397_), .B(new_n729_), .C1(new_n490_), .C2(new_n512_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n733_), .A2(new_n650_), .A3(new_n669_), .A4(new_n706_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G99gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(KEYINPUT109), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT51), .B1(new_n743_), .B2(KEYINPUT109), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n743_), .A2(KEYINPUT108), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(G1338gat));
  NAND4_X1  g547(.A1(new_n733_), .A2(new_n256_), .A3(new_n669_), .A4(new_n706_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G106gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G106gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n256_), .A2(new_n203_), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n751_), .A2(new_n752_), .B1(new_n729_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g554(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n617_), .B2(new_n448_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n580_), .A2(new_n449_), .A3(new_n616_), .A4(new_n756_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n428_), .A2(new_n429_), .A3(new_n438_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n430_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT114), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n427_), .A2(new_n765_), .A3(new_n439_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n766_), .A3(new_n434_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n444_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n445_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT115), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n772_), .A3(new_n445_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n612_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n608_), .A2(new_n448_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT111), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n591_), .B2(KEYINPUT112), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n592_), .A2(new_n596_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n586_), .B1(new_n782_), .B2(new_n584_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n591_), .A2(KEYINPUT112), .A3(new_n779_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(KEYINPUT113), .A3(KEYINPUT56), .A4(new_n610_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n608_), .A2(new_n788_), .A3(new_n448_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n778_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n591_), .A2(KEYINPUT112), .A3(new_n779_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n792_), .A2(new_n780_), .A3(new_n783_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(new_n611_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n776_), .B1(new_n790_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n761_), .B1(new_n798_), .B2(new_n624_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n797_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n778_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n775_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(KEYINPUT57), .A3(new_n625_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n774_), .A2(new_n608_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n774_), .A2(new_n608_), .A3(KEYINPUT117), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n807_), .A2(new_n808_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n579_), .B(new_n804_), .C1(new_n809_), .C2(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n808_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT117), .B1(new_n774_), .B2(new_n608_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n793_), .A2(new_n791_), .A3(new_n611_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n610_), .ZN(new_n816_));
  OAI22_X1  g615(.A1(new_n813_), .A2(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n804_), .B1(new_n819_), .B2(new_n579_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n799_), .B(new_n803_), .C1(new_n812_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n626_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n807_), .A2(new_n808_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n794_), .A2(new_n796_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT58), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT118), .B1(new_n826_), .B2(new_n666_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n811_), .A3(new_n810_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT119), .A3(new_n803_), .A4(new_n799_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT120), .B(new_n760_), .C1(new_n823_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n821_), .A2(new_n822_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n480_), .A3(new_n829_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n760_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n831_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n830_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n642_), .A2(new_n256_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n350_), .A3(new_n650_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n448_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n828_), .A2(new_n799_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n828_), .A2(KEYINPUT121), .A3(new_n799_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n803_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n760_), .B1(new_n847_), .B2(new_n480_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(KEYINPUT59), .A3(new_n838_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n840_), .B2(KEYINPUT59), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n449_), .A2(KEYINPUT122), .ZN(new_n851_));
  MUX2_X1   g650(.A(KEYINPUT122), .B(new_n851_), .S(G113gat), .Z(new_n852_));
  AOI21_X1  g651(.A(new_n842_), .B1(new_n850_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n616_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n841_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n616_), .B(new_n849_), .C1(new_n840_), .C2(KEYINPUT59), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n841_), .A2(new_n859_), .A3(new_n626_), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n480_), .B(new_n849_), .C1(new_n840_), .C2(KEYINPUT59), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n841_), .B2(new_n624_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT123), .B(G134gat), .Z(new_n864_));
  NOR2_X1   g663(.A1(new_n666_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n850_), .B2(new_n865_), .ZN(G1343gat));
  NAND3_X1  g665(.A1(new_n256_), .A2(new_n350_), .A3(new_n397_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n830_), .A2(new_n835_), .A3(new_n642_), .A4(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n448_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n627_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n626_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n868_), .A2(new_n876_), .A3(new_n624_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n868_), .A2(new_n579_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n876_), .ZN(G1347gat));
  OR3_X1    g678(.A1(new_n655_), .A2(new_n641_), .A3(new_n374_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n848_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n448_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT62), .B1(new_n882_), .B2(KEYINPUT22), .ZN(new_n883_));
  OAI21_X1  g682(.A(G169gat), .B1(new_n882_), .B2(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(G169gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n883_), .ZN(G1348gat));
  AOI21_X1  g686(.A(G176gat), .B1(new_n881_), .B2(new_n627_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n836_), .A2(KEYINPUT124), .A3(new_n255_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT124), .B1(new_n836_), .B2(new_n255_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n641_), .A2(new_n374_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n892_), .A2(G176gat), .A3(new_n627_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n891_), .B2(new_n893_), .ZN(G1349gat));
  AND3_X1   g693(.A1(new_n881_), .A2(new_n301_), .A3(new_n626_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n626_), .B(new_n892_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n272_), .ZN(G1350gat));
  NAND4_X1  g696(.A1(new_n881_), .A2(new_n275_), .A3(new_n280_), .A4(new_n624_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n848_), .A2(new_n666_), .A3(new_n880_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n274_), .B2(new_n899_), .ZN(G1351gat));
  NAND2_X1  g699(.A1(new_n833_), .A2(new_n834_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT120), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n833_), .A2(new_n831_), .A3(new_n834_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n642_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(new_n903_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT125), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n902_), .A2(new_n908_), .A3(new_n903_), .A4(new_n905_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G197gat), .B1(new_n910_), .B2(new_n448_), .ZN(new_n911_));
  INV_X1    g710(.A(G197gat), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n912_), .B(new_n449_), .C1(new_n907_), .C2(new_n909_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n627_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(G204gat), .ZN(new_n916_));
  INV_X1    g715(.A(G204gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n910_), .A2(new_n917_), .A3(new_n627_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1353gat));
  NOR3_X1   g718(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n480_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n922_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n908_), .B1(new_n836_), .B2(new_n905_), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n830_), .A2(new_n835_), .A3(KEYINPUT125), .A4(new_n904_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n923_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(new_n926_), .A3(new_n921_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n910_), .A2(new_n934_), .A3(new_n624_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n666_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(new_n936_), .ZN(G1355gat));
endmodule


