//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n993_, new_n994_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1020_, new_n1021_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT10), .B(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT64), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n205_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n217_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n217_), .A2(new_n215_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n213_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n225_), .B1(new_n205_), .B2(new_n230_), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n214_), .A2(new_n223_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233_));
  INV_X1    g032(.A(new_n229_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(KEYINPUT66), .A3(new_n229_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .A3(new_n225_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  XOR2_X1   g041(.A(G71gat), .B(G78gat), .Z(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n232_), .A2(new_n240_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n211_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT64), .B1(new_n209_), .B2(new_n210_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n213_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n223_), .A3(new_n238_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n231_), .A2(new_n224_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n240_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n247_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n202_), .B1(new_n249_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n255_), .B2(new_n247_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n249_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI211_X1 g060(.A(new_n258_), .B(KEYINPUT12), .C1(new_n255_), .C2(new_n247_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n257_), .B1(new_n263_), .B2(new_n202_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G176gat), .B(G204gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT69), .ZN(new_n266_));
  XOR2_X1   g065(.A(G120gat), .B(G148gat), .Z(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  OR3_X1    g069(.A1(new_n264_), .A2(KEYINPUT70), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n248_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT12), .B1(new_n272_), .B2(new_n258_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n260_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n273_), .A2(new_n202_), .A3(new_n249_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n257_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n270_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n270_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT70), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n271_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT13), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n271_), .A2(KEYINPUT13), .A3(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT71), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G29gat), .B(G36gat), .Z(new_n289_));
  XOR2_X1   g088(.A(G43gat), .B(G50gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G29gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G43gat), .B(G50gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT15), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G1gat), .A2(G8gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n297_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G15gat), .ZN(new_n304_));
  INV_X1    g103(.A(G22gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G15gat), .A2(G22gat), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(KEYINPUT14), .B2(new_n301_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n300_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n303_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n303_), .B2(new_n309_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n296_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n308_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n309_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n315_), .B1(new_n316_), .B2(new_n302_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n317_), .A2(new_n310_), .B1(new_n294_), .B2(new_n291_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n311_), .A2(new_n295_), .A3(new_n312_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(new_n318_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n295_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n310_), .A3(new_n317_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n319_), .A2(new_n327_), .A3(KEYINPUT75), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n320_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n322_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AOI211_X1 g130(.A(KEYINPUT76), .B(new_n320_), .C1(new_n325_), .C2(new_n328_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n321_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G141gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G169gat), .B(G197gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(KEYINPUT77), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  OAI221_X1 g137(.A(new_n321_), .B1(KEYINPUT77), .B2(new_n336_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT18), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT90), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT90), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  INV_X1    g157(.A(G176gat), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n355_), .A2(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT23), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G183gat), .ZN(new_n366_));
  INV_X1    g165(.A(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n365_), .A2(KEYINPUT91), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT91), .B1(new_n365_), .B2(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n364_), .A3(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n361_), .A2(KEYINPUT23), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT80), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(G169gat), .B2(G176gat), .ZN(new_n379_));
  INV_X1    g178(.A(G169gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n359_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n366_), .A2(KEYINPUT25), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G183gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT26), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G190gat), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n376_), .A2(new_n382_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n371_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G204gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT84), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G204gat), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT21), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(G197gat), .B2(G204gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n398_), .A2(KEYINPUT85), .A3(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G218gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G211gat), .ZN(new_n407_));
  INV_X1    g206(.A(G211gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G218gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G197gat), .A2(G204gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(G204gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n397_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT21), .B1(new_n410_), .B2(KEYINPUT87), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G211gat), .B(G218gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n414_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n405_), .A2(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n352_), .B1(new_n392_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n389_), .A2(KEYINPUT78), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT25), .B(G183gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G190gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT78), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n426_), .A2(new_n365_), .A3(new_n382_), .A4(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n373_), .A2(new_n375_), .A3(new_n368_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(G176gat), .B1(new_n433_), .B2(KEYINPUT22), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT22), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n354_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n425_), .B1(new_n423_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n397_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n415_), .B1(new_n441_), .B2(new_n411_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n398_), .A2(KEYINPUT85), .A3(new_n400_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT85), .B1(new_n398_), .B2(new_n400_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n442_), .B(new_n418_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n421_), .A2(new_n422_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n431_), .A2(new_n438_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(KEYINPUT92), .A3(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n424_), .A2(KEYINPUT97), .B1(new_n440_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n391_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n351_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n376_), .A2(new_n455_), .A3(new_n382_), .A4(new_n389_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n381_), .A2(KEYINPUT24), .A3(new_n353_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n377_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n389_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n373_), .A2(new_n375_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT89), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n371_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n447_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n352_), .B1(new_n423_), .B2(new_n439_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n464_), .A2(new_n351_), .A3(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT98), .B(new_n348_), .C1(new_n454_), .C2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT98), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n440_), .A2(new_n449_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n447_), .C2(new_n391_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n453_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n466_), .B1(new_n471_), .B2(new_n350_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n468_), .B1(new_n472_), .B2(new_n347_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G1gat), .B(G29gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT96), .B(G85gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT0), .B(G57gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NAND2_X1  g278(.A1(G225gat), .A2(G233gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(G127gat), .B(G134gat), .Z(new_n481_));
  XOR2_X1   g280(.A(G113gat), .B(G120gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G141gat), .A2(G148gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G141gat), .A2(G148gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT2), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G155gat), .A2(G162gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT82), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G155gat), .A3(G162gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G155gat), .A2(G162gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT83), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n504_), .A3(new_n501_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n494_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n488_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n485_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n500_), .B1(new_n499_), .B2(KEYINPUT1), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT1), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n496_), .A2(new_n498_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n484_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(KEYINPUT1), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n501_), .A3(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n508_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n504_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n518_));
  AOI211_X1 g317(.A(KEYINPUT83), .B(new_n500_), .C1(new_n496_), .C2(new_n498_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n493_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n520_), .A3(new_n483_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(KEYINPUT4), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n514_), .A2(KEYINPUT94), .A3(KEYINPUT4), .A4(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n514_), .B2(KEYINPUT4), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n517_), .A2(new_n520_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT4), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n529_), .A2(KEYINPUT95), .A3(new_n530_), .A4(new_n484_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n480_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n514_), .A2(new_n521_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n480_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n479_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n538_));
  INV_X1    g337(.A(new_n479_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n528_), .A2(new_n531_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n539_), .B(new_n540_), .C1(new_n542_), .C2(new_n480_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n533_), .A2(new_n536_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT99), .A3(new_n539_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n351_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n351_), .A2(KEYINPUT20), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n363_), .B1(G183gat), .B2(G190gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n368_), .B1(new_n549_), .B2(new_n374_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n365_), .A2(KEYINPUT91), .A3(new_n368_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n456_), .A2(new_n461_), .B1(new_n554_), .B2(new_n360_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n548_), .B1(new_n555_), .B2(new_n423_), .ZN(new_n556_));
  AOI221_X4 g355(.A(new_n425_), .B1(new_n431_), .B2(new_n438_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT92), .B1(new_n447_), .B2(new_n448_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT93), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n556_), .B(new_n561_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n547_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n347_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n474_), .A2(new_n544_), .A3(new_n546_), .A4(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n562_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n547_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n346_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AOI211_X1 g367(.A(new_n547_), .B(new_n345_), .C1(new_n560_), .C2(new_n562_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT33), .B(new_n479_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n537_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n542_), .A2(new_n480_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n479_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n565_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G227gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n304_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G71gat), .B(G99gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(G43gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(G43gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT30), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n582_), .A2(G43gat), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n583_), .ZN(new_n589_));
  AND4_X1   g388(.A1(new_n438_), .A2(new_n431_), .A3(new_n586_), .A4(new_n589_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n438_), .A2(new_n431_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n581_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n448_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n431_), .A2(new_n586_), .A3(new_n438_), .A4(new_n589_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n580_), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT31), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT31), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n592_), .A2(new_n593_), .A3(new_n600_), .A4(new_n597_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n599_), .A2(new_n484_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n484_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G228gat), .A2(G233gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n529_), .A2(KEYINPUT29), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n607_), .B2(new_n447_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n606_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n610_), .A2(new_n423_), .A3(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(KEYINPUT88), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n517_), .A2(new_n520_), .A3(new_n609_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT28), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT28), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n517_), .A2(new_n520_), .A3(new_n618_), .A4(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G22gat), .B(G50gat), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G78gat), .B(G106gat), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT88), .B1(new_n608_), .B2(new_n612_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n625_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n615_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n625_), .A2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n626_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n625_), .A2(new_n628_), .A3(new_n627_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n614_), .A3(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n605_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n578_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n562_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n561_), .B1(new_n469_), .B2(new_n556_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n567_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n345_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n563_), .A2(new_n346_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT27), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n345_), .B1(new_n454_), .B2(new_n466_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n563_), .B2(new_n346_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n644_), .A2(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n544_), .A2(new_n546_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n604_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n602_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n603_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n631_), .A2(new_n635_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n648_), .B(new_n649_), .C1(new_n650_), .C2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n341_), .B1(new_n638_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT34), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT35), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n296_), .A2(new_n255_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(KEYINPUT72), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n326_), .B2(new_n255_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G190gat), .B(G218gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT73), .ZN(new_n664_));
  XOR2_X1   g463(.A(G134gat), .B(G162gat), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n661_), .A2(new_n662_), .B1(KEYINPUT36), .B2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n657_), .A2(KEYINPUT35), .ZN(new_n668_));
  OAI221_X1 g467(.A(new_n659_), .B1(new_n326_), .B2(new_n255_), .C1(new_n660_), .C2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n666_), .A2(KEYINPUT36), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n667_), .B(new_n669_), .C1(KEYINPUT36), .C2(new_n666_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT37), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(KEYINPUT37), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(G231gat), .A2(G233gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n247_), .B(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(new_n313_), .ZN(new_n681_));
  XOR2_X1   g480(.A(G127gat), .B(G155gat), .Z(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT16), .ZN(new_n683_));
  XNOR2_X1  g482(.A(G183gat), .B(G211gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT17), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n685_), .B(KEYINPUT17), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n681_), .B2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n678_), .A2(new_n691_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n288_), .A2(new_n655_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n649_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT100), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n649_), .A2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n693_), .A2(new_n298_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT101), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n693_), .A2(new_n702_), .A3(new_n298_), .A4(new_n699_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(KEYINPUT38), .A3(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT102), .Z(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT38), .B1(new_n701_), .B2(new_n703_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n286_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(new_n341_), .A3(new_n691_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n674_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n638_), .B2(new_n654_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n298_), .B1(new_n711_), .B2(new_n694_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n706_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n705_), .A2(new_n713_), .ZN(G1324gat));
  INV_X1    g513(.A(new_n648_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n299_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT39), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n693_), .A2(new_n299_), .A3(new_n715_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g519(.A(new_n304_), .B1(new_n711_), .B2(new_n604_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT41), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n693_), .A2(new_n304_), .A3(new_n604_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n631_), .A2(new_n635_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n305_), .B1(new_n711_), .B2(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT42), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n693_), .A2(new_n305_), .A3(new_n725_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1327gat));
  INV_X1    g528(.A(new_n691_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n674_), .A2(new_n730_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n655_), .A2(new_n286_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G29gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n694_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n286_), .A2(new_n340_), .A3(new_n691_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n650_), .A2(new_n653_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n644_), .A2(new_n645_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n647_), .A2(new_n646_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n649_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n636_), .B1(new_n565_), .B2(new_n577_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n678_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT43), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n638_), .A2(new_n654_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n678_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n737_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n736_), .B1(new_n749_), .B2(KEYINPUT44), .ZN(new_n750_));
  INV_X1    g549(.A(new_n737_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n747_), .B1(new_n746_), .B2(new_n678_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n678_), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT43), .B(new_n753_), .C1(new_n638_), .C2(new_n654_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(KEYINPUT103), .A3(new_n756_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n750_), .A2(new_n757_), .B1(KEYINPUT44), .B2(new_n749_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n699_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n735_), .B1(new_n759_), .B2(G29gat), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT104), .B(new_n733_), .C1(new_n758_), .C2(new_n699_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n734_), .B1(new_n760_), .B2(new_n761_), .ZN(G1328gat));
  INV_X1    g561(.A(G36gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n732_), .A2(new_n763_), .A3(new_n715_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT45), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT44), .B(new_n751_), .C1(new_n752_), .C2(new_n754_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n715_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n749_), .A2(new_n736_), .A3(KEYINPUT44), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT103), .B1(new_n755_), .B2(new_n756_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT105), .B1(new_n771_), .B2(G36gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n767_), .B1(new_n750_), .B2(new_n757_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n763_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n765_), .B1(new_n772_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT46), .B(new_n765_), .C1(new_n772_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1329gat));
  NAND3_X1  g579(.A1(new_n758_), .A2(G43gat), .A3(new_n604_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n732_), .A2(new_n604_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(G43gat), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g583(.A(G50gat), .B1(new_n732_), .B2(new_n725_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n725_), .A2(G50gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n758_), .B2(new_n786_), .ZN(G1331gat));
  NOR3_X1   g586(.A1(new_n288_), .A2(new_n340_), .A3(new_n691_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n710_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G57gat), .B1(new_n789_), .B2(new_n649_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n746_), .A2(new_n341_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT107), .Z(new_n792_));
  NAND2_X1  g591(.A1(new_n707_), .A2(new_n692_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT106), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT108), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n698_), .A2(G57gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n790_), .B1(new_n796_), .B2(new_n797_), .ZN(G1332gat));
  OAI21_X1  g597(.A(G64gat), .B1(new_n789_), .B2(new_n648_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT48), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n648_), .A2(G64gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n796_), .B2(new_n801_), .ZN(G1333gat));
  OAI21_X1  g601(.A(G71gat), .B1(new_n789_), .B2(new_n605_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT49), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n605_), .A2(G71gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n796_), .B2(new_n805_), .ZN(G1334gat));
  INV_X1    g605(.A(new_n725_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G78gat), .B1(new_n789_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT50), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n807_), .A2(G78gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n796_), .B2(new_n810_), .ZN(G1335gat));
  AND2_X1   g610(.A1(new_n287_), .A2(new_n731_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n792_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G85gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n699_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n745_), .A2(new_n748_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n286_), .A2(new_n340_), .A3(new_n730_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818_), .B2(new_n649_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(G1336gat));
  INV_X1    g619(.A(G92gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n821_), .A3(new_n715_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G92gat), .B1(new_n818_), .B2(new_n648_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1337gat));
  NAND3_X1  g623(.A1(new_n813_), .A2(new_n604_), .A3(new_n212_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G99gat), .B1(new_n818_), .B2(new_n605_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(KEYINPUT109), .A3(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829_));
  INV_X1    g628(.A(new_n818_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT111), .A3(new_n725_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G106gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT111), .B1(new_n830_), .B2(new_n725_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n833_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n831_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n807_), .A2(G106gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n792_), .A2(new_n812_), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT110), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT53), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n834_), .A2(new_n836_), .A3(new_n839_), .A4(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1339gat));
  NOR3_X1   g643(.A1(new_n678_), .A2(new_n340_), .A3(new_n691_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n286_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(KEYINPUT54), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(KEYINPUT54), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n336_), .B(new_n321_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n330_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n336_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n314_), .A2(new_n319_), .A3(new_n330_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n851_), .B2(new_n336_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n271_), .A2(new_n281_), .A3(new_n850_), .A4(new_n856_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n338_), .A2(new_n339_), .B1(new_n264_), .B2(new_n270_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n860_));
  NAND2_X1  g659(.A1(new_n275_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n261_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n862_), .A2(KEYINPUT55), .A3(new_n202_), .A4(new_n274_), .ZN(new_n863_));
  OAI211_X1 g662(.A(G230gat), .B(G233gat), .C1(new_n261_), .C2(new_n262_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n859_), .B1(new_n865_), .B2(new_n278_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n858_), .B1(new_n866_), .B2(KEYINPUT56), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n859_), .B(new_n868_), .C1(new_n865_), .C2(new_n278_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n857_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n674_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(KEYINPUT57), .A3(new_n674_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n865_), .A2(new_n278_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT56), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n865_), .A2(new_n868_), .A3(new_n278_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n856_), .A2(new_n280_), .A3(new_n850_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n877_), .A2(KEYINPUT58), .A3(new_n878_), .A4(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n678_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n856_), .A2(new_n280_), .A3(new_n850_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n876_), .B2(KEYINPUT56), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT58), .B1(new_n883_), .B2(new_n878_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n875_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(KEYINPUT116), .A3(new_n678_), .A4(new_n880_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n873_), .A2(new_n874_), .A3(new_n885_), .A4(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n730_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n885_), .A2(new_n889_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n870_), .A2(KEYINPUT57), .A3(new_n674_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n872_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n870_), .B2(new_n674_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n897_), .A3(KEYINPUT117), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n849_), .B1(new_n892_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n699_), .A2(new_n648_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(KEYINPUT118), .A3(new_n650_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903_));
  INV_X1    g702(.A(new_n650_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n900_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT59), .B1(new_n899_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n906_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909_));
  INV_X1    g708(.A(new_n849_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n876_), .A2(KEYINPUT113), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n868_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n866_), .A2(KEYINPUT56), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n913_), .A3(new_n858_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n709_), .B1(new_n914_), .B2(new_n857_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n874_), .B1(new_n915_), .B2(new_n895_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n881_), .A2(new_n884_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n691_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n908_), .A2(new_n909_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n907_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G113gat), .B1(new_n921_), .B2(new_n341_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n885_), .A2(new_n889_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n891_), .B1(new_n916_), .B2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n898_), .A2(new_n924_), .A3(new_n691_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n910_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n926_), .A2(new_n927_), .A3(new_n908_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT119), .B1(new_n899_), .B2(new_n906_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n341_), .A2(G113gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n922_), .B1(new_n930_), .B2(new_n931_), .ZN(G1340gat));
  OAI21_X1  g731(.A(G120gat), .B1(new_n921_), .B2(new_n288_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934_));
  AOI21_X1  g733(.A(G120gat), .B1(new_n707_), .B2(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT120), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n934_), .B2(G120gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n928_), .A2(new_n929_), .A3(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n939_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n933_), .B1(new_n940_), .B2(new_n941_), .ZN(G1341gat));
  OAI21_X1  g741(.A(G127gat), .B1(new_n921_), .B2(new_n691_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n691_), .A2(G127gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n930_), .B2(new_n944_), .ZN(G1342gat));
  INV_X1    g744(.A(new_n921_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n678_), .A2(G134gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT122), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n928_), .A2(new_n929_), .A3(new_n709_), .ZN(new_n949_));
  INV_X1    g748(.A(G134gat), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n946_), .A2(new_n948_), .B1(new_n949_), .B2(new_n950_), .ZN(G1343gat));
  INV_X1    g750(.A(new_n653_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n899_), .A2(new_n952_), .A3(new_n900_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n340_), .ZN(new_n954_));
  XOR2_X1   g753(.A(KEYINPUT123), .B(G141gat), .Z(new_n955_));
  XNOR2_X1  g754(.A(new_n954_), .B(new_n955_), .ZN(G1344gat));
  NAND2_X1  g755(.A1(new_n953_), .A2(new_n287_), .ZN(new_n957_));
  XOR2_X1   g756(.A(KEYINPUT124), .B(G148gat), .Z(new_n958_));
  XNOR2_X1  g757(.A(new_n957_), .B(new_n958_), .ZN(G1345gat));
  AOI21_X1  g758(.A(new_n952_), .B1(new_n925_), .B2(new_n910_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n960_), .A2(new_n730_), .A3(new_n901_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(KEYINPUT125), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n953_), .A2(new_n963_), .A3(new_n730_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(KEYINPUT61), .B(G155gat), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n967_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n962_), .A2(new_n964_), .A3(new_n966_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1346gat));
  INV_X1    g769(.A(new_n953_), .ZN(new_n971_));
  OR3_X1    g770(.A1(new_n971_), .A2(G162gat), .A3(new_n674_), .ZN(new_n972_));
  OAI21_X1  g771(.A(G162gat), .B1(new_n971_), .B2(new_n753_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(G1347gat));
  NAND3_X1  g773(.A1(new_n698_), .A2(new_n604_), .A3(new_n715_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n975_), .A2(new_n725_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n919_), .A2(new_n976_), .ZN(new_n977_));
  INV_X1    g776(.A(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n380_), .B1(new_n978_), .B2(new_n340_), .ZN(new_n979_));
  OR2_X1    g778(.A1(new_n979_), .A2(KEYINPUT62), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n978_), .A2(new_n340_), .A3(new_n358_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n979_), .A2(KEYINPUT62), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n980_), .A2(new_n981_), .A3(new_n982_), .ZN(G1348gat));
  AOI21_X1  g782(.A(G176gat), .B1(new_n978_), .B2(new_n707_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n899_), .A2(new_n725_), .ZN(new_n985_));
  NOR3_X1   g784(.A1(new_n288_), .A2(new_n359_), .A3(new_n975_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n984_), .B1(new_n985_), .B2(new_n986_), .ZN(G1349gat));
  NOR3_X1   g786(.A1(new_n977_), .A2(new_n427_), .A3(new_n691_), .ZN(new_n988_));
  NOR4_X1   g787(.A1(new_n899_), .A2(new_n725_), .A3(new_n691_), .A4(new_n975_), .ZN(new_n989_));
  OR2_X1    g788(.A1(new_n989_), .A2(KEYINPUT126), .ZN(new_n990_));
  AOI21_X1  g789(.A(G183gat), .B1(new_n989_), .B2(KEYINPUT126), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n988_), .B1(new_n990_), .B2(new_n991_), .ZN(G1350gat));
  OAI21_X1  g791(.A(G190gat), .B1(new_n977_), .B2(new_n753_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n709_), .A2(new_n428_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n977_), .B2(new_n994_), .ZN(G1351gat));
  NOR2_X1   g794(.A1(new_n694_), .A2(new_n648_), .ZN(new_n996_));
  NAND3_X1  g795(.A1(new_n926_), .A2(new_n653_), .A3(new_n996_), .ZN(new_n997_));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n997_), .A2(new_n998_), .ZN(new_n999_));
  NAND3_X1  g798(.A1(new_n960_), .A2(KEYINPUT127), .A3(new_n996_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n999_), .A2(new_n1000_), .ZN(new_n1001_));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001_), .B2(new_n340_), .ZN(new_n1002_));
  AOI211_X1 g801(.A(new_n397_), .B(new_n341_), .C1(new_n999_), .C2(new_n1000_), .ZN(new_n1003_));
  NOR2_X1   g802(.A1(new_n1002_), .A2(new_n1003_), .ZN(G1352gat));
  INV_X1    g803(.A(new_n413_), .ZN(new_n1005_));
  AOI21_X1  g804(.A(KEYINPUT127), .B1(new_n960_), .B2(new_n996_), .ZN(new_n1006_));
  INV_X1    g805(.A(new_n996_), .ZN(new_n1007_));
  NOR4_X1   g806(.A1(new_n899_), .A2(new_n998_), .A3(new_n952_), .A4(new_n1007_), .ZN(new_n1008_));
  OAI211_X1 g807(.A(new_n1005_), .B(new_n287_), .C1(new_n1006_), .C2(new_n1008_), .ZN(new_n1009_));
  AOI21_X1  g808(.A(new_n288_), .B1(new_n999_), .B2(new_n1000_), .ZN(new_n1010_));
  OAI21_X1  g809(.A(new_n1009_), .B1(new_n1010_), .B2(G204gat), .ZN(new_n1011_));
  INV_X1    g810(.A(new_n1011_), .ZN(G1353gat));
  NOR2_X1   g811(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1013_));
  INV_X1    g812(.A(new_n1013_), .ZN(new_n1014_));
  AOI21_X1  g813(.A(new_n691_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1015_));
  AOI21_X1  g814(.A(new_n1014_), .B1(new_n1001_), .B2(new_n1015_), .ZN(new_n1016_));
  INV_X1    g815(.A(new_n1015_), .ZN(new_n1017_));
  AOI211_X1 g816(.A(new_n1013_), .B(new_n1017_), .C1(new_n999_), .C2(new_n1000_), .ZN(new_n1018_));
  NOR2_X1   g817(.A1(new_n1016_), .A2(new_n1018_), .ZN(G1354gat));
  NAND3_X1  g818(.A1(new_n1001_), .A2(new_n406_), .A3(new_n709_), .ZN(new_n1020_));
  AOI21_X1  g819(.A(new_n753_), .B1(new_n999_), .B2(new_n1000_), .ZN(new_n1021_));
  OAI21_X1  g820(.A(new_n1020_), .B1(new_n406_), .B2(new_n1021_), .ZN(G1355gat));
endmodule


