//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n565_, new_n566_, new_n567_, new_n568_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G29gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT87), .B(G127gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G134gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n207_), .B(new_n208_), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT96), .ZN(new_n210_));
  AND2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G141gat), .ZN(new_n216_));
  INV_X1    g015(.A(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n218_), .B(KEYINPUT3), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n219_), .B(KEYINPUT2), .Z(new_n225_));
  OAI21_X1  g024(.A(new_n213_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n207_), .B(new_n208_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT96), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n210_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT97), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n227_), .A2(new_n228_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(KEYINPUT97), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT98), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n235_), .B2(KEYINPUT4), .ZN(new_n240_));
  INV_X1    g039(.A(new_n236_), .ZN(new_n241_));
  OAI221_X1 g040(.A(new_n205_), .B1(new_n235_), .B2(new_n237_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G169gat), .ZN(new_n243_));
  INV_X1    g042(.A(G176gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(KEYINPUT24), .A3(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(KEYINPUT24), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT23), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT26), .B(G190gat), .Z(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT25), .B(G183gat), .Z(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n246_), .A2(KEYINPUT93), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n258_), .B2(new_n244_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n256_), .B(new_n257_), .C1(KEYINPUT93), .C2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G197gat), .B(G204gat), .Z(new_n262_));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT21), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n264_), .B(new_n265_), .C1(KEYINPUT21), .C2(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n261_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT94), .ZN(new_n271_));
  INV_X1    g070(.A(new_n253_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT83), .B(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(KEYINPUT25), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n252_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n259_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n251_), .B1(new_n274_), .B2(G190gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n259_), .A2(new_n279_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n284_), .B2(new_n268_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n271_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n261_), .A2(new_n269_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT95), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n268_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(KEYINPUT95), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n288_), .A2(KEYINPUT20), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n292_), .B(KEYINPUT92), .Z(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT19), .Z(new_n294_));
  MUX2_X1   g093(.A(new_n286_), .B(new_n291_), .S(new_n294_), .Z(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT18), .B(G64gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G92gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n295_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT99), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n240_), .A2(new_n302_), .A3(new_n237_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n205_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n235_), .A2(new_n241_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n302_), .B1(new_n240_), .B2(new_n237_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(KEYINPUT100), .A3(KEYINPUT33), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT33), .B1(new_n307_), .B2(KEYINPUT100), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n242_), .B(new_n301_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT101), .ZN(new_n312_));
  INV_X1    g111(.A(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n308_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT101), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n242_), .A4(new_n301_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT103), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(new_n205_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(new_n307_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n307_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n287_), .A2(KEYINPUT20), .A3(new_n289_), .ZN(new_n322_));
  MUX2_X1   g121(.A(new_n322_), .B(new_n286_), .S(new_n294_), .Z(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT32), .A3(new_n299_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT32), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n295_), .B1(new_n325_), .B2(new_n300_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT102), .Z(new_n327_));
  NAND4_X1  g126(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .A4(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n312_), .A2(new_n316_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n268_), .B1(new_n227_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G228gat), .ZN(new_n332_));
  INV_X1    g131(.A(G233gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT91), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G78gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n227_), .A2(new_n330_), .ZN(new_n338_));
  INV_X1    g137(.A(G106gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n337_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT91), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n341_), .B(new_n342_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n228_), .B(KEYINPUT31), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n284_), .B(KEYINPUT30), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G71gat), .B(G99gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G15gat), .B(G43gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n356_), .B(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n329_), .A2(new_n351_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n351_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n347_), .A2(new_n350_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n320_), .A2(new_n321_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n301_), .A2(KEYINPUT27), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT104), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n295_), .A2(new_n299_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n323_), .A2(new_n300_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT27), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n368_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n363_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G85gat), .B(G92gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G99gat), .A2(G106gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT6), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G99gat), .A3(G106gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT7), .ZN(new_n387_));
  INV_X1    g186(.A(G99gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n339_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT67), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n391_), .A2(new_n387_), .A3(new_n388_), .A4(new_n339_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT66), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT66), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n390_), .A2(new_n392_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n386_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT8), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT70), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n390_), .A2(new_n392_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n381_), .B1(G99gat), .B2(G106gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n379_), .A2(KEYINPUT6), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT69), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n394_), .A2(new_n396_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n401_), .A2(new_n404_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n378_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT8), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n380_), .A2(new_n382_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n397_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n400_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n408_), .A2(KEYINPUT9), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT10), .B(G99gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT64), .B(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(KEYINPUT9), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(G85gat), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n417_), .A2(new_n420_), .A3(new_n424_), .A4(new_n412_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n416_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G57gat), .B(G64gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(KEYINPUT11), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(KEYINPUT11), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G78gat), .ZN(new_n430_));
  OR3_X1    g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n430_), .A3(KEYINPUT11), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n426_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT12), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n416_), .A2(new_n425_), .A3(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G230gat), .A2(G233gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n426_), .A2(KEYINPUT12), .A3(new_n434_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT72), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n435_), .A2(new_n444_), .A3(new_n438_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n439_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n426_), .A2(KEYINPUT71), .A3(new_n434_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n443_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G120gat), .B(G148gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(G204gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT5), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(new_n244_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(KEYINPUT73), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n443_), .A2(new_n448_), .A3(new_n453_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n449_), .A2(new_n453_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n460_), .A2(KEYINPUT13), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(KEYINPUT13), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G15gat), .B(G22gat), .Z(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT80), .B(G1gat), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G8gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n466_), .B2(KEYINPUT14), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G1gat), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n468_), .A2(G8gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(G8gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  INV_X1    g272(.A(G43gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G50gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n471_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n476_), .B(KEYINPUT15), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n472_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(new_n243_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G197gat), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT82), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n487_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n463_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n377_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT34), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT75), .Z(new_n499_));
  AND2_X1   g298(.A1(new_n484_), .A2(new_n426_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n416_), .A2(new_n425_), .A3(new_n478_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n496_), .A2(new_n497_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n500_), .B1(new_n503_), .B2(KEYINPUT76), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(KEYINPUT76), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n499_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n501_), .B(new_n502_), .C1(KEYINPUT77), .C2(new_n499_), .ZN(new_n507_));
  AOI211_X1 g306(.A(new_n507_), .B(new_n500_), .C1(KEYINPUT77), .C2(new_n499_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G190gat), .B(G218gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G134gat), .ZN(new_n510_));
  INV_X1    g309(.A(G162gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OR4_X1    g312(.A1(KEYINPUT36), .A2(new_n506_), .A3(new_n508_), .A4(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n512_), .B(KEYINPUT36), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT79), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT106), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT106), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G231gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n433_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n471_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT16), .B(G183gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G211gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G127gat), .B(G155gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n529_), .A2(new_n530_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n525_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n531_), .B2(new_n525_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n522_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n494_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(G1gat), .B1(new_n538_), .B2(new_n369_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n517_), .B2(KEYINPUT78), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n518_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n514_), .B(new_n517_), .C1(KEYINPUT78), .C2(new_n540_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n463_), .A2(new_n535_), .A3(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT81), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n492_), .B1(new_n545_), .B2(KEYINPUT81), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n377_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n369_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(KEYINPUT105), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(KEYINPUT105), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(new_n465_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT38), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n539_), .A2(new_n555_), .ZN(G1324gat));
  INV_X1    g355(.A(G8gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n375_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n537_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g363(.A(G15gat), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n537_), .B2(new_n364_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT41), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n548_), .A2(new_n565_), .A3(new_n364_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(G1326gat));
  INV_X1    g368(.A(G22gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n548_), .A2(new_n570_), .A3(new_n366_), .ZN(new_n571_));
  OAI21_X1  g370(.A(G22gat), .B1(new_n538_), .B2(new_n351_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(KEYINPUT42), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(KEYINPUT42), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n571_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT108), .ZN(G1327gat));
  INV_X1    g375(.A(KEYINPUT43), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n377_), .B2(new_n544_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n377_), .A2(new_n577_), .A3(new_n544_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n535_), .A3(new_n493_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT44), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n581_), .A2(KEYINPUT44), .A3(new_n535_), .A4(new_n493_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n552_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(G29gat), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n521_), .A2(new_n534_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT109), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n494_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT110), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n494_), .A2(KEYINPUT110), .A3(new_n591_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n369_), .A2(G29gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT111), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n589_), .B1(new_n597_), .B2(new_n599_), .ZN(G1328gat));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n558_), .A3(new_n585_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G36gat), .ZN(new_n602_));
  INV_X1    g401(.A(G36gat), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n594_), .A2(new_n603_), .A3(new_n558_), .A4(new_n595_), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT46), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(G1329gat));
  NAND3_X1  g408(.A1(new_n594_), .A2(new_n364_), .A3(new_n595_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT113), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n474_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n610_), .B2(new_n474_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AND4_X1   g413(.A1(G43gat), .A2(new_n584_), .A3(new_n364_), .A4(new_n585_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n614_), .A2(new_n615_), .A3(KEYINPUT47), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT47), .B1(new_n614_), .B2(new_n615_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1330gat));
  AOI21_X1  g417(.A(G50gat), .B1(new_n596_), .B2(new_n366_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n586_), .A2(new_n366_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n620_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g420(.A(new_n463_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n492_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n363_), .B2(new_n376_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n535_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G57gat), .B1(new_n628_), .B2(new_n587_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n626_), .A2(new_n536_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n549_), .A2(G57gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(G1332gat));
  INV_X1    g431(.A(G64gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n630_), .B2(new_n558_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT48), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n633_), .A3(new_n558_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1333gat));
  INV_X1    g436(.A(G71gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n630_), .B2(new_n364_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT114), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT49), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n628_), .A2(new_n638_), .A3(new_n364_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1334gat));
  AOI21_X1  g442(.A(new_n336_), .B1(new_n630_), .B2(new_n366_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT115), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT50), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n628_), .A2(new_n336_), .A3(new_n366_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1335gat));
  AND2_X1   g447(.A1(new_n626_), .A2(new_n591_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G85gat), .B1(new_n649_), .B2(new_n587_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n544_), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT43), .B(new_n651_), .C1(new_n363_), .C2(new_n376_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n535_), .B(new_n624_), .C1(new_n578_), .C2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(G85gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n650_), .B1(new_n655_), .B2(new_n549_), .ZN(G1336gat));
  AOI21_X1  g455(.A(G92gat), .B1(new_n649_), .B2(new_n558_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n423_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n375_), .B1(new_n658_), .B2(new_n421_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n654_), .B2(new_n659_), .ZN(G1337gat));
  OAI21_X1  g459(.A(G99gat), .B1(new_n653_), .B2(new_n362_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n649_), .A2(new_n418_), .A3(new_n364_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT51), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n661_), .A2(new_n662_), .B1(KEYINPUT116), .B2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT116), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1338gat));
  AOI21_X1  g465(.A(new_n625_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT117), .A3(new_n535_), .A4(new_n366_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT117), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n653_), .B2(new_n351_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n670_), .A3(G106gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT52), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT52), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n668_), .A2(new_n670_), .A3(new_n673_), .A4(G106gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n649_), .A2(new_n419_), .A3(new_n366_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT53), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT53), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1339gat));
  INV_X1    g480(.A(KEYINPUT121), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n492_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT55), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n442_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT119), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT12), .B1(new_n426_), .B2(new_n434_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n436_), .B(new_n433_), .C1(new_n416_), .C2(new_n425_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n689_), .B2(new_n438_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n438_), .ZN(new_n691_));
  NOR4_X1   g490(.A1(new_n687_), .A2(new_n688_), .A3(new_n691_), .A4(KEYINPUT119), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n685_), .B1(new_n693_), .B2(new_n446_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT72), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n689_), .B2(new_n440_), .ZN(new_n696_));
  AND4_X1   g495(.A1(new_n695_), .A2(new_n437_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n684_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT118), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT118), .B(new_n684_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n453_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(KEYINPUT56), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT56), .B1(new_n702_), .B2(new_n703_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n683_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT120), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n485_), .A2(new_n479_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n482_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n477_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n490_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n487_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n490_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n460_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT120), .B(new_n683_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n708_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n521_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT57), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(KEYINPUT57), .A3(new_n521_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n458_), .B(new_n714_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT58), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n544_), .A3(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n721_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n535_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n492_), .B(new_n627_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT54), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n682_), .B1(new_n728_), .B2(new_n732_), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT121), .B(new_n731_), .C1(new_n727_), .C2(new_n535_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n552_), .A2(new_n558_), .A3(new_n365_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n733_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G113gat), .B1(new_n737_), .B2(new_n623_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n731_), .B1(new_n727_), .B2(new_n535_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n736_), .A2(new_n739_), .A3(KEYINPUT59), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT122), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT59), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n737_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n728_), .A2(new_n732_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT121), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n739_), .A2(new_n682_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n735_), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n740_), .B1(new_n743_), .B2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n623_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n738_), .B1(new_n750_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g550(.A(KEYINPUT123), .ZN(new_n752_));
  INV_X1    g551(.A(G120gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n749_), .B2(new_n463_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n737_), .B(new_n755_), .C1(KEYINPUT60), .C2(new_n753_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n752_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n740_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n737_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT122), .B1(new_n747_), .B2(KEYINPUT59), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n463_), .B(new_n759_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G120gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(KEYINPUT123), .A3(new_n756_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n758_), .A2(new_n764_), .ZN(G1341gat));
  AOI21_X1  g564(.A(G127gat), .B1(new_n737_), .B2(new_n534_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n749_), .A2(G127gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(new_n534_), .ZN(G1342gat));
  NAND2_X1  g567(.A1(new_n544_), .A2(G134gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT124), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n759_), .B(new_n770_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n771_));
  INV_X1    g570(.A(G134gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n747_), .B2(new_n521_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT125), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT125), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(new_n776_), .A3(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1343gat));
  NOR3_X1   g577(.A1(new_n733_), .A2(new_n734_), .A3(new_n367_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n552_), .A2(new_n558_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(new_n492_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(new_n216_), .ZN(G1344gat));
  NOR2_X1   g582(.A1(new_n781_), .A2(new_n622_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(new_n217_), .ZN(G1345gat));
  NOR2_X1   g584(.A1(new_n781_), .A2(new_n535_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT61), .B(G155gat), .Z(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(G1346gat));
  NOR3_X1   g587(.A1(new_n781_), .A2(new_n511_), .A3(new_n651_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(new_n522_), .A3(new_n780_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n511_), .B2(new_n790_), .ZN(G1347gat));
  NAND3_X1  g590(.A1(new_n552_), .A2(new_n364_), .A3(new_n558_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n739_), .A2(new_n366_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n623_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G169gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT62), .ZN(new_n796_));
  INV_X1    g595(.A(new_n258_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n794_), .ZN(G1348gat));
  AOI21_X1  g597(.A(G176gat), .B1(new_n793_), .B2(new_n463_), .ZN(new_n799_));
  OR4_X1    g598(.A1(new_n366_), .A2(new_n733_), .A3(new_n734_), .A4(new_n792_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n244_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n801_), .B2(new_n463_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT126), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1349gat));
  AND3_X1   g603(.A1(new_n793_), .A2(new_n534_), .A3(new_n254_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n800_), .A2(new_n535_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n273_), .ZN(G1350gat));
  NAND2_X1  g606(.A1(new_n522_), .A2(new_n272_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT127), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n793_), .A2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n793_), .A2(new_n544_), .ZN(new_n811_));
  INV_X1    g610(.A(G190gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(G1351gat));
  NAND2_X1  g612(.A1(new_n779_), .A2(new_n558_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n549_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n623_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n463_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n534_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT63), .B(G211gat), .Z(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(new_n822_), .ZN(G1354gat));
  AOI21_X1  g622(.A(G218gat), .B1(new_n815_), .B2(new_n522_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n815_), .A2(G218gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n544_), .B2(new_n825_), .ZN(G1355gat));
endmodule


