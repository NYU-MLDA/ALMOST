//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT25), .B(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT79), .B1(new_n209_), .B2(KEYINPUT26), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n208_), .B(new_n210_), .C1(new_n211_), .C2(KEYINPUT79), .ZN(new_n212_));
  OR3_X1    g011(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n212_), .A2(new_n203_), .A3(new_n213_), .A4(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n207_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G43gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G71gat), .B(G99gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT30), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G227gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G15gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n223_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n221_), .B(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT80), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  INV_X1    g028(.A(G113gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G120gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(G113gat), .ZN(new_n233_));
  INV_X1    g032(.A(G120gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT31), .Z(new_n237_));
  OR2_X1    g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(KEYINPUT80), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G197gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT85), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(KEYINPUT86), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n245_), .B(KEYINPUT87), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n249_), .B(new_n250_), .C1(KEYINPUT21), .C2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n250_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT89), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT84), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT2), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT82), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT3), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT3), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n268_), .B(KEYINPUT83), .C1(new_n271_), .C2(new_n272_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n266_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n264_), .A2(new_n278_), .A3(KEYINPUT1), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n264_), .B2(KEYINPUT1), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n279_), .A2(new_n263_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n269_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n282_), .A2(new_n267_), .A3(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n277_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n242_), .B1(new_n262_), .B2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n258_), .A2(new_n242_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G78gat), .B(G106gat), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n257_), .B(KEYINPUT89), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(new_n287_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n299_), .A2(new_n242_), .B1(new_n291_), .B2(new_n290_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n294_), .ZN(new_n301_));
  OR3_X1    g100(.A1(new_n277_), .A2(KEYINPUT29), .A3(new_n284_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT28), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(KEYINPUT28), .ZN(new_n304_));
  XOR2_X1   g103(.A(G22gat), .B(G50gat), .Z(new_n305_));
  AND3_X1   g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AND4_X1   g107(.A1(KEYINPUT90), .A2(new_n296_), .A3(new_n301_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n300_), .B2(new_n294_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n311_), .A2(new_n308_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT93), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n232_), .A2(new_n235_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n236_), .A2(KEYINPUT93), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n285_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n236_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(new_n314_), .C1(new_n284_), .C2(new_n277_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n285_), .A2(new_n318_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n320_), .A2(KEYINPUT4), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n323_), .B1(new_n326_), .B2(new_n322_), .ZN(new_n327_));
  XOR2_X1   g126(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G57gat), .B(G85gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(KEYINPUT33), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT96), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n327_), .A2(new_n332_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT33), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT97), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n254_), .A2(new_n256_), .A3(new_n207_), .A4(new_n219_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n211_), .A2(new_n208_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n339_), .A2(new_n218_), .A3(new_n203_), .A4(new_n213_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT92), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT92), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n342_), .A2(new_n343_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT20), .B(new_n338_), .C1(new_n344_), .C2(new_n258_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT91), .Z(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT19), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n258_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n257_), .A2(new_n220_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n351_), .A2(KEYINPUT20), .A3(new_n348_), .A4(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G64gat), .ZN(new_n357_));
  INV_X1    g156(.A(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n359_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n337_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n326_), .A2(KEYINPUT98), .A3(new_n322_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n332_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n326_), .A2(new_n322_), .ZN(new_n368_));
  OAI221_X1 g167(.A(new_n367_), .B1(KEYINPUT98), .B2(new_n368_), .C1(new_n322_), .C2(new_n321_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n335_), .A2(KEYINPUT97), .A3(new_n336_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n334_), .A2(new_n364_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n345_), .A2(new_n349_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT100), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n207_), .A2(new_n340_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT99), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n297_), .C2(new_n375_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n352_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n372_), .B1(new_n380_), .B2(new_n349_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT101), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT101), .ZN(new_n384_));
  INV_X1    g183(.A(new_n382_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n352_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n375_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n377_), .B1(new_n262_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n388_), .B2(KEYINPUT100), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n348_), .B1(new_n389_), .B2(new_n378_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n384_), .B(new_n385_), .C1(new_n390_), .C2(new_n372_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n327_), .A2(new_n332_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n335_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n354_), .A2(new_n382_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n383_), .A2(new_n391_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n313_), .B1(new_n371_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n393_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n350_), .A2(new_n353_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n359_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n401_), .B2(new_n361_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT102), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT102), .B(new_n398_), .C1(new_n401_), .C2(new_n361_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT27), .B(new_n360_), .C1(new_n381_), .C2(new_n359_), .ZN(new_n407_));
  AND4_X1   g206(.A1(new_n397_), .A2(new_n313_), .A3(new_n406_), .A4(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n241_), .B1(new_n396_), .B2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n406_), .A2(new_n407_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n313_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n393_), .A2(new_n241_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G230gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G85gat), .B(G92gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT9), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G99gat), .A2(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT6), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(G99gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(KEYINPUT10), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(KEYINPUT10), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n425_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G85gat), .ZN(new_n430_));
  OR3_X1    g229(.A1(new_n430_), .A2(new_n358_), .A3(KEYINPUT9), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n419_), .A2(new_n424_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI211_X1 g235(.A(KEYINPUT8), .B(new_n417_), .C1(new_n436_), .C2(new_n424_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n426_), .A3(new_n425_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n422_), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n420_), .A2(KEYINPUT6), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n433_), .B(new_n440_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n438_), .B1(new_n443_), .B2(new_n418_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n432_), .B1(new_n437_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT64), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n447_), .B(new_n432_), .C1(new_n437_), .C2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  XOR2_X1   g250(.A(G71gat), .B(G78gat), .Z(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n443_), .A2(new_n418_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT8), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n443_), .A2(new_n438_), .A3(new_n418_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n429_), .A2(new_n424_), .A3(new_n431_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n459_), .A2(new_n460_), .B1(new_n419_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n449_), .A2(new_n457_), .B1(new_n463_), .B2(KEYINPUT12), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n446_), .A2(new_n448_), .A3(new_n456_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n466_));
  AND3_X1   g265(.A1(new_n465_), .A2(KEYINPUT67), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT67), .B1(new_n465_), .B2(new_n466_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n416_), .B(new_n464_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n449_), .A2(new_n457_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT65), .A3(new_n465_), .ZN(new_n472_));
  OR3_X1    g271(.A1(new_n449_), .A2(KEYINPUT65), .A3(new_n457_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n416_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G120gat), .B(G148gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT5), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G176gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(new_n246_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n476_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n469_), .A2(new_n475_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(new_n481_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT69), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT13), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(KEYINPUT68), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n469_), .A2(new_n475_), .A3(new_n470_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n481_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n485_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n476_), .A2(new_n477_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT69), .B1(new_n496_), .B2(new_n481_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT13), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  INV_X1    g300(.A(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT74), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n504_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G1gat), .B(G8gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G29gat), .B(G36gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(G43gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(G43gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G50gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(G50gat), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT77), .ZN(new_n523_));
  INV_X1    g322(.A(new_n512_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525_));
  INV_X1    g324(.A(new_n519_), .ZN(new_n526_));
  AOI21_X1  g325(.A(G50gat), .B1(new_n514_), .B2(new_n515_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT15), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n523_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n520_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n523_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  MUX2_X1   g335(.A(new_n532_), .B(new_n534_), .S(new_n536_), .Z(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT78), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n216_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n244_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n537_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n500_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n415_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n459_), .A2(new_n460_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n447_), .B1(new_n546_), .B2(new_n432_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n448_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n521_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n530_), .A2(new_n445_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n549_), .A2(new_n552_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n520_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n462_), .B1(new_n529_), .B2(new_n528_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT35), .B(new_n551_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT70), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G134gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G162gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n565_), .A2(KEYINPUT71), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n565_), .A2(KEYINPUT71), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n558_), .B(new_n555_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n559_), .A2(KEYINPUT72), .A3(new_n565_), .A4(new_n566_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n574_), .A2(new_n575_), .A3(KEYINPUT37), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n574_), .B2(KEYINPUT37), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n567_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT37), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n512_), .B(new_n457_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT75), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n582_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G183gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(G211gat), .Z(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n585_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n590_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n581_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT76), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n545_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n501_), .A3(new_n393_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT38), .ZN(new_n603_));
  INV_X1    g402(.A(new_n579_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n596_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n545_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n397_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(G1324gat));
  OAI21_X1  g407(.A(G8gat), .B1(new_n606_), .B2(new_n410_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT39), .ZN(new_n610_));
  INV_X1    g409(.A(new_n410_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n601_), .A2(new_n502_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n606_), .B2(new_n241_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n241_), .A2(G15gat), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n600_), .B2(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n606_), .B2(new_n411_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n411_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n600_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT104), .ZN(G1327gat));
  INV_X1    g423(.A(new_n581_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n415_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT43), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT43), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n415_), .A2(new_n628_), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(KEYINPUT44), .A3(new_n544_), .A4(new_n596_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n415_), .B2(new_n625_), .ZN(new_n632_));
  AOI211_X1 g431(.A(KEYINPUT43), .B(new_n581_), .C1(new_n409_), .C2(new_n414_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n544_), .B(new_n596_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G29gat), .B1(new_n637_), .B2(new_n397_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n597_), .A2(new_n579_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n545_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n397_), .A2(G29gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT105), .Z(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n640_), .B2(new_n642_), .ZN(G1328gat));
  OAI21_X1  g442(.A(KEYINPUT106), .B1(new_n637_), .B2(new_n410_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n631_), .A2(new_n636_), .A3(new_n645_), .A4(new_n611_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(G36gat), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n640_), .A2(G36gat), .A3(new_n410_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n647_), .B(new_n650_), .C1(KEYINPUT108), .C2(KEYINPUT46), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  INV_X1    g454(.A(new_n241_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n631_), .A2(new_n636_), .A3(G43gat), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(G43gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n640_), .B2(new_n241_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT109), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(KEYINPUT47), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1330gat));
  OAI21_X1  g467(.A(G50gat), .B1(new_n637_), .B2(new_n411_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n313_), .A2(new_n517_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n640_), .B2(new_n670_), .ZN(G1331gat));
  NOR2_X1   g470(.A1(new_n499_), .A2(new_n542_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n605_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(G57gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT110), .B1(new_n397_), .B2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n676_), .A2(KEYINPUT110), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n678_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(new_n393_), .A3(new_n599_), .A4(new_n674_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n681_), .B2(new_n677_), .ZN(G1332gat));
  OAI21_X1  g481(.A(G64gat), .B1(new_n675_), .B2(new_n410_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT48), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n674_), .A2(new_n599_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n410_), .A2(G64gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(G1333gat));
  OAI21_X1  g486(.A(G71gat), .B1(new_n675_), .B2(new_n241_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT49), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n241_), .A2(G71gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n685_), .B2(new_n690_), .ZN(G1334gat));
  OR3_X1    g490(.A1(new_n685_), .A2(G78gat), .A3(new_n411_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G78gat), .B1(new_n675_), .B2(new_n411_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT111), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(G78gat), .C1(new_n675_), .C2(new_n411_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n694_), .A2(KEYINPUT50), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT50), .B1(new_n694_), .B2(new_n696_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n692_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT112), .Z(G1335gat));
  OAI211_X1 g499(.A(new_n596_), .B(new_n672_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n701_), .A2(new_n430_), .A3(new_n397_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n674_), .A2(new_n639_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT113), .Z(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n393_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n705_), .B2(new_n430_), .ZN(G1336gat));
  NOR3_X1   g505(.A1(new_n701_), .A2(new_n358_), .A3(new_n410_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n611_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(new_n358_), .ZN(G1337gat));
  OAI211_X1 g508(.A(new_n704_), .B(new_n656_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT115), .ZN(new_n711_));
  OAI21_X1  g510(.A(G99gat), .B1(new_n701_), .B2(new_n241_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(KEYINPUT114), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n710_), .B(new_n713_), .C1(KEYINPUT114), .C2(new_n712_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(G1338gat));
  AOI21_X1  g515(.A(new_n673_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n717_), .A2(KEYINPUT117), .A3(new_n313_), .A4(new_n596_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT117), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n701_), .B2(new_n411_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n720_), .A3(G106gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT52), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n718_), .A2(new_n720_), .A3(new_n723_), .A4(G106gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n704_), .A2(new_n425_), .A3(new_n313_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n729_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  NOR3_X1   g530(.A1(new_n495_), .A2(new_n497_), .A3(KEYINPUT13), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n487_), .B1(new_n486_), .B2(new_n492_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n543_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT118), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n598_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT119), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n734_), .B2(new_n598_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n542_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n596_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT118), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n737_), .B1(new_n741_), .B2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT119), .B1(new_n744_), .B2(KEYINPUT54), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n736_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n464_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n752_), .A2(KEYINPUT120), .A3(new_n474_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT120), .B1(new_n752_), .B2(new_n474_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n469_), .B(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT121), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n752_), .A2(new_n474_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n752_), .A2(KEYINPUT120), .A3(new_n474_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n469_), .B(KEYINPUT55), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT121), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n758_), .A2(new_n481_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT56), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n758_), .A2(new_n769_), .A3(new_n766_), .A4(new_n481_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n768_), .A2(new_n542_), .A3(new_n494_), .A4(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT122), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT122), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n523_), .A2(new_n536_), .A3(new_n531_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n534_), .A2(new_n536_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n541_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n774_), .A2(new_n776_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT123), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n772_), .A2(new_n773_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n751_), .B1(new_n781_), .B2(new_n604_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n768_), .A2(new_n494_), .A3(new_n770_), .A4(new_n777_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n784_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n581_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n768_), .A2(new_n770_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n542_), .A4(new_n494_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n771_), .A2(KEYINPUT122), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n778_), .B(KEYINPUT123), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n579_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n782_), .A2(new_n788_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n750_), .B1(new_n796_), .B2(new_n596_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n412_), .A2(new_n393_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n797_), .A2(new_n241_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n542_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n750_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n579_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT57), .B1(new_n794_), .B2(new_n579_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n787_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n804_), .B2(new_n597_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT59), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n798_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n656_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n797_), .B2(KEYINPUT124), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n799_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n543_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n800_), .B1(new_n814_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g614(.A(new_n234_), .B1(new_n499_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n799_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n234_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n499_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n234_), .ZN(G1341gat));
  AOI21_X1  g618(.A(G127gat), .B1(new_n799_), .B2(new_n597_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n596_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g621(.A(G134gat), .B1(new_n799_), .B2(new_n604_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n581_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g624(.A1(new_n797_), .A2(new_n411_), .A3(new_n611_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n397_), .A2(new_n656_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n542_), .A3(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n500_), .A3(new_n827_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n597_), .A3(new_n827_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT61), .B(G155gat), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1346gat));
  NOR2_X1   g633(.A1(new_n611_), .A2(new_n411_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n805_), .A2(new_n835_), .A3(new_n604_), .A4(new_n827_), .ZN(new_n836_));
  INV_X1    g635(.A(G162gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT125), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n840_), .A3(new_n837_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n826_), .A2(new_n827_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n581_), .A2(new_n837_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n839_), .A2(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(G1347gat));
  NAND2_X1  g643(.A1(new_n411_), .A2(new_n413_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n805_), .A2(new_n611_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT126), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n796_), .A2(new_n596_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n410_), .B1(new_n849_), .B2(new_n801_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT126), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n846_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT22), .B(G169gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n848_), .A2(new_n542_), .A3(new_n852_), .A4(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n542_), .A3(new_n846_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(G169gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n855_), .B2(G169gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(G1348gat));
  NOR3_X1   g658(.A1(new_n847_), .A2(new_n217_), .A3(new_n499_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n848_), .A2(new_n500_), .A3(new_n852_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n217_), .ZN(G1349gat));
  NOR2_X1   g661(.A1(new_n847_), .A2(new_n596_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(G183gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n851_), .B1(new_n850_), .B2(new_n846_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n797_), .A2(KEYINPUT126), .A3(new_n410_), .A4(new_n845_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n596_), .A2(new_n208_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n867_), .B2(new_n868_), .ZN(G1350gat));
  NAND4_X1  g668(.A1(new_n848_), .A2(new_n211_), .A3(new_n852_), .A4(new_n604_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n865_), .A2(new_n866_), .A3(new_n581_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n209_), .ZN(G1351gat));
  NOR3_X1   g671(.A1(new_n411_), .A2(new_n393_), .A3(new_n656_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n850_), .A2(new_n542_), .A3(new_n873_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n874_), .A2(KEYINPUT127), .A3(new_n244_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT127), .B1(new_n874_), .B2(new_n244_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n244_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(G1352gat));
  NAND2_X1  g677(.A1(new_n805_), .A2(new_n611_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n873_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n879_), .A2(new_n499_), .A3(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n246_), .ZN(G1353gat));
  NAND3_X1  g681(.A1(new_n850_), .A2(new_n597_), .A3(new_n873_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  AND2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n883_), .B2(new_n884_), .ZN(G1354gat));
  NOR2_X1   g686(.A1(new_n879_), .A2(new_n880_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G218gat), .B1(new_n888_), .B2(new_n604_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n625_), .A2(G218gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n888_), .B2(new_n890_), .ZN(G1355gat));
endmodule


