//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n205_));
  OR2_X1    g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n202_), .A2(new_n203_), .A3(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT10), .B(G99gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n209_), .B(new_n212_), .C1(G106gat), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT7), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT66), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n222_), .A2(new_n224_), .A3(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n206_), .A2(new_n202_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n215_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n215_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n212_), .B2(new_n222_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n214_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n242_), .B(new_n214_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n235_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G230gat), .ZN(new_n250_));
  INV_X1    g049(.A(G233gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n244_), .A2(new_n245_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n252_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G120gat), .B(G148gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(new_n256_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n256_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n252_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(KEYINPUT68), .B(new_n263_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT13), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n270_), .A2(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT13), .B1(new_n268_), .B2(new_n269_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT69), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT78), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G29gat), .A2(G36gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G29gat), .A2(G36gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(G43gat), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(G29gat), .A2(G36gat), .ZN(new_n285_));
  INV_X1    g084(.A(G43gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n281_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G50gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(new_n287_), .A3(G50gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n302_), .A2(KEYINPUT77), .A3(new_n303_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT15), .ZN(new_n311_));
  INV_X1    g110(.A(new_n291_), .ZN(new_n312_));
  AOI21_X1  g111(.A(G50gat), .B1(new_n284_), .B2(new_n287_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n290_), .A2(KEYINPUT15), .A3(new_n291_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n300_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n307_), .A3(new_n302_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G141gat), .ZN(new_n319_));
  INV_X1    g118(.A(G169gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G197gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n310_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n310_), .B2(new_n318_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n280_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT78), .A3(new_n325_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n279_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G57gat), .B(G85gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  NAND3_X1  g144(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  OR3_X1    g148(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G141gat), .ZN(new_n358_));
  INV_X1    g157(.A(G148gat), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n352_), .A2(KEYINPUT1), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n357_), .A2(new_n344_), .A3(new_n346_), .A4(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G127gat), .A2(G134gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G127gat), .A2(G134gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(G113gat), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G127gat), .ZN(new_n366_));
  INV_X1    g165(.A(G134gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G113gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n362_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n370_), .A3(G120gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n370_), .ZN(new_n372_));
  INV_X1    g171(.A(G120gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n355_), .A2(new_n361_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT91), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n355_), .A2(new_n361_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n365_), .A2(new_n370_), .A3(G120gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(G120gat), .B1(new_n365_), .B2(new_n370_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(KEYINPUT81), .A3(new_n371_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n376_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .A4(KEYINPUT91), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(KEYINPUT4), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n344_), .A2(new_n346_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n392_), .A2(new_n360_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n379_), .A2(new_n380_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n386_), .B1(new_n388_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n389_), .B1(new_n396_), .B2(KEYINPUT4), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n341_), .B(new_n387_), .C1(new_n397_), .C2(new_n385_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n385_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n403_), .B2(new_n389_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n404_), .A2(KEYINPUT33), .A3(new_n341_), .A4(new_n387_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n384_), .A2(new_n401_), .A3(new_n386_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(new_n340_), .C1(new_n397_), .C2(new_n401_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n400_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT18), .B(G64gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT19), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT20), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G190gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT87), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n419_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G183gat), .A2(G190gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT23), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n320_), .A2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT24), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(KEYINPUT24), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n426_), .A2(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(G183gat), .B2(G190gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n427_), .A2(KEYINPUT23), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n436_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n432_), .ZN(new_n441_));
  OR2_X1    g240(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443_));
  NAND2_X1  g242(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT88), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(G176gat), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n441_), .A2(new_n449_), .A3(KEYINPUT89), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451_));
  INV_X1    g250(.A(new_n432_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n428_), .B2(new_n436_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT88), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n443_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n429_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n435_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(G211gat), .A2(G218gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G211gat), .A2(G218gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT21), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G197gat), .B(G204gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT21), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n465_), .A3(new_n460_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n463_), .A3(KEYINPUT21), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n417_), .B1(new_n458_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n429_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT79), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n429_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n472_), .A2(new_n440_), .A3(new_n432_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n422_), .A2(new_n418_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n476_), .A2(new_n428_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n475_), .A2(KEYINPUT80), .A3(new_n477_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n469_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n416_), .B1(new_n470_), .B2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n426_), .A2(new_n434_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(new_n469_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT89), .B1(new_n441_), .B2(new_n449_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n453_), .A2(new_n456_), .A3(new_n451_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n417_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n475_), .A2(KEYINPUT80), .A3(new_n477_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT80), .B1(new_n475_), .B2(new_n477_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n469_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n416_), .A3(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n413_), .B1(new_n484_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n497_), .B2(new_n482_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n483_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n415_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n490_), .A2(new_n416_), .A3(new_n493_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n412_), .A3(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n495_), .A2(new_n496_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n496_), .B1(new_n495_), .B2(new_n502_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n408_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT95), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n435_), .B(new_n482_), .C1(new_n441_), .C2(new_n449_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n493_), .A2(new_n511_), .A3(KEYINPUT20), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n415_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n470_), .A2(new_n416_), .A3(new_n483_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n507_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n510_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT96), .B(new_n507_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n509_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n404_), .A2(new_n341_), .A3(new_n387_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n341_), .B1(new_n404_), .B2(new_n387_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT97), .B1(new_n519_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(new_n516_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT96), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n515_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n404_), .A2(new_n387_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n340_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n398_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n527_), .A2(new_n530_), .A3(new_n531_), .A4(new_n509_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n506_), .A2(new_n523_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n381_), .A2(new_n382_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT31), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G227gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(G15gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G43gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT30), .B1(new_n491_), .B2(new_n492_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n480_), .A2(new_n543_), .A3(new_n481_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G71gat), .B(G99gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n542_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n541_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT30), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n543_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n545_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n542_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n540_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT82), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT82), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n536_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT84), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G228gat), .A2(G233gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n469_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT84), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(new_n469_), .C1(new_n393_), .C2(new_n560_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G78gat), .B(G106gat), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT85), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n393_), .A2(new_n560_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G22gat), .B(G50gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT28), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n575_), .B(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n570_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT86), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT86), .A4(new_n578_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n557_), .B1(new_n549_), .B2(new_n554_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n535_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n559_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n533_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT27), .B1(new_n495_), .B2(new_n502_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n515_), .A2(new_n413_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(new_n502_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n594_), .B2(KEYINPUT27), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n549_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n535_), .B1(new_n596_), .B2(new_n588_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n556_), .A2(new_n536_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n587_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n587_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n522_), .B(new_n595_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n591_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n235_), .A2(new_n316_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n293_), .B(new_n214_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n606_), .A2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n603_), .A2(new_n609_), .A3(new_n613_), .A4(new_n608_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(KEYINPUT72), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(KEYINPUT36), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n607_), .B(new_n606_), .C1(new_n603_), .C2(new_n609_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n614_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT36), .B(new_n620_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n621_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n612_), .A2(KEYINPUT72), .A3(new_n626_), .A4(new_n614_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n628_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT37), .B1(new_n628_), .B2(KEYINPUT73), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT75), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(G183gat), .B(G211gat), .Z(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n637_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n639_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n633_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n643_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(KEYINPUT17), .A3(new_n641_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n242_), .B(new_n300_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n243_), .A2(new_n300_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n301_), .A2(new_n242_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n648_), .A3(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n644_), .B(new_n646_), .C1(new_n649_), .C2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n642_), .A2(new_n633_), .A3(new_n643_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n647_), .A2(new_n648_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n651_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(G231gat), .A3(G233gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n653_), .A2(new_n658_), .A3(KEYINPUT76), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT76), .B1(new_n653_), .B2(new_n658_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n632_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n333_), .A2(new_n602_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT98), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n295_), .A3(new_n530_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT38), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n582_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n668_), .B1(new_n559_), .B2(new_n589_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n597_), .A2(new_n598_), .A3(new_n587_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n530_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n671_), .A2(new_n595_), .B1(new_n533_), .B2(new_n590_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n653_), .A2(new_n658_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n672_), .A2(new_n628_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n333_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT99), .Z(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n530_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n667_), .B1(new_n295_), .B2(new_n677_), .ZN(G1324gat));
  INV_X1    g477(.A(new_n595_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n674_), .A2(new_n333_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(G8gat), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT39), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n682_), .A2(new_n686_), .A3(G8gat), .A4(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n665_), .A2(new_n296_), .A3(new_n679_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT102), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1325gat));
  NOR2_X1   g495(.A1(new_n559_), .A2(new_n589_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n665_), .A2(new_n538_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n676_), .A2(new_n698_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n700_), .B2(G15gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(G1326gat));
  INV_X1    g502(.A(G22gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n665_), .A2(new_n704_), .A3(new_n587_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n676_), .A2(new_n587_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G22gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT42), .B(new_n704_), .C1(new_n676_), .C2(new_n587_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1327gat));
  NAND4_X1  g509(.A1(new_n274_), .A2(new_n278_), .A3(new_n331_), .A4(new_n662_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n628_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n711_), .A2(new_n672_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n530_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT103), .B1(new_n629_), .B2(new_n630_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n628_), .A2(KEYINPUT73), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT37), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n628_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n672_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n602_), .A2(new_n725_), .A3(new_n632_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n711_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n715_), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n591_), .B2(new_n601_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n632_), .A2(new_n725_), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n729_), .A2(new_n725_), .B1(new_n672_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n711_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(KEYINPUT104), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n728_), .A2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(G29gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n727_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n522_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n714_), .B1(new_n737_), .B2(new_n741_), .ZN(G1328gat));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n595_), .B1(new_n728_), .B2(new_n735_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n740_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n713_), .A2(new_n743_), .A3(new_n679_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT45), .Z(new_n749_));
  OR3_X1    g548(.A1(new_n746_), .A2(new_n747_), .A3(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1329gat));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT105), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n754_));
  AND4_X1   g553(.A1(KEYINPUT105), .A2(new_n731_), .A3(KEYINPUT44), .A4(new_n732_), .ZN(new_n755_));
  OAI211_X1 g554(.A(G43gat), .B(new_n698_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT104), .B1(new_n733_), .B2(new_n734_), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n715_), .B(KEYINPUT44), .C1(new_n731_), .C2(new_n732_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n713_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n286_), .B1(new_n761_), .B2(new_n697_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n286_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(new_n736_), .A3(KEYINPUT106), .A4(new_n698_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT47), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n760_), .A2(new_n764_), .A3(new_n767_), .A4(new_n762_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1330gat));
  NAND3_X1  g568(.A1(new_n745_), .A2(new_n736_), .A3(new_n587_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT107), .B1(new_n770_), .B2(G50gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n587_), .A2(new_n289_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT108), .Z(new_n774_));
  OAI22_X1  g573(.A1(new_n771_), .A2(new_n772_), .B1(new_n761_), .B2(new_n774_), .ZN(G1331gat));
  AND2_X1   g574(.A1(new_n279_), .A2(new_n663_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT109), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT109), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n331_), .A4(new_n672_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G57gat), .B1(new_n779_), .B2(new_n530_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT110), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(KEYINPUT110), .ZN(new_n782_));
  INV_X1    g581(.A(new_n279_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n661_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NOR4_X1   g584(.A1(new_n783_), .A2(new_n672_), .A3(new_n628_), .A4(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n530_), .A2(G57gat), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n781_), .A2(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(G1332gat));
  INV_X1    g587(.A(G64gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n786_), .B2(new_n679_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT48), .Z(new_n791_));
  NAND3_X1  g590(.A1(new_n779_), .A2(new_n789_), .A3(new_n679_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1333gat));
  INV_X1    g592(.A(G71gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n786_), .B2(new_n698_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT49), .Z(new_n796_));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n794_), .A3(new_n698_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1334gat));
  INV_X1    g597(.A(G78gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n786_), .B2(new_n587_), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT50), .Z(new_n801_));
  NAND3_X1  g600(.A1(new_n779_), .A2(new_n799_), .A3(new_n587_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1335gat));
  NAND3_X1  g602(.A1(new_n279_), .A2(new_n332_), .A3(new_n662_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(new_n712_), .A3(new_n672_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT111), .Z(new_n806_));
  AOI21_X1  g605(.A(G85gat), .B1(new_n806_), .B2(new_n530_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n731_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n808_), .A2(new_n804_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT112), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(new_n530_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n807_), .B1(new_n811_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g611(.A(G92gat), .B1(new_n806_), .B2(new_n679_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n810_), .A2(new_n679_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(KEYINPUT51), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(KEYINPUT51), .ZN(new_n818_));
  INV_X1    g617(.A(new_n213_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n806_), .A2(new_n819_), .A3(new_n698_), .ZN(new_n820_));
  OAI21_X1  g619(.A(G99gat), .B1(new_n809_), .B2(new_n697_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n817_), .B(new_n818_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  AND4_X1   g621(.A1(new_n816_), .A2(new_n820_), .A3(KEYINPUT51), .A4(new_n821_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1338gat));
  NAND3_X1  g623(.A1(new_n806_), .A2(new_n217_), .A3(new_n587_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n808_), .A2(new_n668_), .A3(new_n804_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(G106gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(G106gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n825_), .B(new_n832_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  OR3_X1    g633(.A1(new_n265_), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT55), .B1(new_n265_), .B2(KEYINPUT116), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n246_), .A2(KEYINPUT117), .A3(new_n252_), .A4(new_n248_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n835_), .A2(new_n837_), .A3(new_n838_), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n263_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n843_), .A3(new_n263_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n842_), .A2(new_n331_), .A3(new_n262_), .A4(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n306_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n317_), .A2(new_n302_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT118), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n323_), .B(new_n846_), .C1(new_n848_), .C2(new_n307_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n849_), .A2(new_n325_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n269_), .A3(new_n268_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n628_), .B1(new_n845_), .B2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT119), .A3(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n842_), .A2(new_n262_), .A3(new_n850_), .A4(new_n844_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT58), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(new_n857_), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n632_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n853_), .B1(KEYINPUT119), .B2(new_n854_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n673_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT114), .B1(new_n272_), .B2(new_n784_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n784_), .B(KEYINPUT114), .C1(new_n275_), .C2(new_n276_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n866_), .B(new_n631_), .C1(new_n867_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT115), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n277_), .B2(new_n785_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n632_), .B1(new_n873_), .B2(new_n868_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n866_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n631_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT54), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n871_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n865_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n679_), .A2(new_n522_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n669_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n332_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n852_), .B(KEYINPUT57), .ZN(new_n886_));
  INV_X1    g685(.A(new_n862_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n662_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n879_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n883_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n865_), .B2(new_n879_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n331_), .B(new_n892_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n895_));
  MUX2_X1   g694(.A(new_n885_), .B(new_n895_), .S(G113gat), .Z(G1340gat));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G120gat), .B1(new_n897_), .B2(new_n783_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n373_), .B1(new_n783_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n893_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n373_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n901_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n898_), .B1(new_n902_), .B2(new_n903_), .ZN(G1341gat));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n662_), .B(new_n890_), .C1(new_n865_), .C2(new_n879_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(G127gat), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT122), .B(new_n366_), .C1(new_n884_), .C2(new_n662_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n673_), .A2(new_n366_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n892_), .B(new_n909_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n907_), .A2(new_n908_), .A3(new_n910_), .ZN(G1342gat));
  OAI21_X1  g710(.A(new_n367_), .B1(new_n884_), .B2(new_n712_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT123), .B(new_n367_), .C1(new_n884_), .C2(new_n712_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n897_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n631_), .A2(new_n367_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT124), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n914_), .A2(new_n915_), .B1(new_n916_), .B2(new_n918_), .ZN(G1343gat));
  AOI21_X1  g718(.A(new_n670_), .B1(new_n865_), .B2(new_n879_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n920_), .A2(new_n881_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n331_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(G141gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n358_), .A3(new_n331_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1344gat));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n279_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G148gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n921_), .A2(new_n359_), .A3(new_n279_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1345gat));
  NAND3_X1  g728(.A1(new_n920_), .A2(new_n661_), .A3(new_n881_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT61), .B(G155gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1346gat));
  NAND2_X1  g731(.A1(new_n921_), .A2(new_n628_), .ZN(new_n933_));
  INV_X1    g732(.A(G162gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n723_), .A2(new_n934_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n934_), .B1(new_n921_), .B2(new_n935_), .ZN(G1347gat));
  NOR4_X1   g735(.A1(new_n697_), .A2(new_n595_), .A3(new_n530_), .A4(new_n587_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n871_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n939_));
  AOI211_X1 g738(.A(new_n939_), .B(new_n628_), .C1(new_n845_), .C2(new_n851_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n853_), .A2(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n661_), .B1(new_n941_), .B2(new_n862_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n331_), .B(new_n937_), .C1(new_n938_), .C2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(KEYINPUT125), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n889_), .A2(new_n945_), .A3(new_n331_), .A4(new_n937_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n944_), .A2(new_n946_), .A3(G169gat), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT62), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n944_), .A2(new_n946_), .A3(new_n949_), .A4(G169gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n889_), .A2(new_n937_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n331_), .B1(new_n455_), .B2(new_n454_), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n954_), .B(KEYINPUT126), .Z(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n951_), .A2(new_n956_), .ZN(G1348gat));
  AOI21_X1  g756(.A(G176gat), .B1(new_n953_), .B2(new_n279_), .ZN(new_n958_));
  AOI211_X1 g757(.A(new_n429_), .B(new_n783_), .C1(new_n865_), .C2(new_n879_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n958_), .B1(new_n937_), .B2(new_n959_), .ZN(G1349gat));
  INV_X1    g759(.A(G183gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n880_), .A2(new_n661_), .A3(new_n937_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n673_), .ZN(new_n963_));
  AND3_X1   g762(.A1(new_n963_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n961_), .A2(new_n962_), .B1(new_n953_), .B2(new_n964_), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n952_), .B2(new_n631_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n628_), .A2(new_n418_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n952_), .B2(new_n967_), .ZN(G1351gat));
  NOR2_X1   g767(.A1(new_n595_), .A2(new_n530_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n920_), .A2(new_n331_), .A3(new_n969_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g770(.A1(new_n920_), .A2(new_n279_), .A3(new_n969_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(KEYINPUT127), .B(G204gat), .ZN(new_n973_));
  XOR2_X1   g772(.A(new_n972_), .B(new_n973_), .Z(G1353gat));
  NAND3_X1  g773(.A1(new_n920_), .A2(new_n963_), .A3(new_n969_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  AND2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n975_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n978_), .B1(new_n975_), .B2(new_n976_), .ZN(G1354gat));
  AND4_X1   g778(.A1(G218gat), .A2(new_n920_), .A3(new_n632_), .A4(new_n969_), .ZN(new_n980_));
  INV_X1    g779(.A(G218gat), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n920_), .A2(new_n628_), .A3(new_n969_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n980_), .B1(new_n981_), .B2(new_n982_), .ZN(G1355gat));
endmodule


