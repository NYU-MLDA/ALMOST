//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n985_, new_n986_, new_n988_, new_n989_, new_n990_, new_n992_,
    new_n993_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1002_, new_n1003_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n214_), .A2(G85gat), .B1(KEYINPUT9), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n210_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(new_n202_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n203_), .A2(KEYINPUT68), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n220_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n203_), .A2(KEYINPUT68), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n202_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n209_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AOI211_X1 g031(.A(KEYINPUT66), .B(KEYINPUT7), .C1(new_n229_), .C2(new_n209_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n224_), .B(new_n227_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n216_), .A2(KEYINPUT67), .A3(new_n211_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n219_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(new_n216_), .B2(new_n211_), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n212_), .A2(new_n215_), .A3(new_n236_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n219_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n243_), .A2(new_n229_), .A3(new_n209_), .A4(new_n228_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n230_), .A2(new_n231_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n206_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n218_), .B1(new_n239_), .B2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G71gat), .B(G78gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(KEYINPUT11), .B2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n253_), .B(new_n218_), .C1(new_n239_), .C2(new_n247_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G230gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT64), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT69), .ZN(new_n261_));
  NAND2_X1  g060(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n255_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n248_), .A2(new_n254_), .A3(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n263_), .A2(new_n264_), .A3(new_n256_), .A4(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n257_), .A2(new_n268_), .A3(new_n259_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n261_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G176gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n261_), .A2(new_n267_), .A3(new_n269_), .A4(new_n275_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n277_), .A2(KEYINPUT13), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT13), .B1(new_n277_), .B2(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G29gat), .B(G36gat), .ZN(new_n283_));
  INV_X1    g082(.A(G43gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT71), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n283_), .B(G43gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n289_), .A3(G50gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(G50gat), .B1(new_n286_), .B2(new_n289_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G8gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT14), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n294_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT73), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n301_), .B(new_n294_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n304_), .A3(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n293_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT15), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n286_), .A2(new_n289_), .ZN(new_n314_));
  INV_X1    g113(.A(G50gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT15), .A3(new_n290_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n308_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n311_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n308_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n290_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n310_), .B1(new_n322_), .B2(new_n309_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G113gat), .B(G141gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G197gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT76), .B(G169gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI22_X1  g127(.A1(new_n319_), .A2(new_n323_), .B1(KEYINPUT75), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n309_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n310_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n328_), .A2(KEYINPUT75), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n291_), .A2(new_n292_), .A3(new_n312_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT15), .B1(new_n316_), .B2(new_n290_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n320_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n282_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT0), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G57gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G85gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G134gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G127gat), .ZN(new_n349_));
  INV_X1    g148(.A(G127gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G134gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G120gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G113gat), .ZN(new_n354_));
  INV_X1    g153(.A(G113gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G120gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n349_), .A2(new_n351_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT86), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT85), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G141gat), .A3(G148gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT2), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373_));
  INV_X1    g172(.A(G141gat), .ZN(new_n374_));
  INV_X1    g173(.A(G148gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n364_), .B(new_n367_), .C1(new_n372_), .C2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n362_), .A2(KEYINPUT1), .B1(new_n374_), .B2(new_n375_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n365_), .A2(new_n382_), .A3(new_n361_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n369_), .A2(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n360_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n372_), .A2(new_n379_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n367_), .A2(new_n364_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n360_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n380_), .A2(new_n385_), .A3(new_n360_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(KEYINPUT97), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n380_), .A2(new_n399_), .A3(new_n385_), .A4(new_n360_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n391_), .B1(new_n401_), .B2(KEYINPUT4), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n390_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n347_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n387_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n405_), .B(new_n346_), .C1(new_n406_), .C2(new_n391_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT27), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT19), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  AND3_X1   g218(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G169gat), .ZN(new_n423_));
  INV_X1    g222(.A(G176gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT24), .A3(new_n426_), .ZN(new_n427_));
  OR3_X1    g226(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT95), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT26), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(G190gat), .ZN(new_n432_));
  INV_X1    g231(.A(G190gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT26), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n430_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT25), .B(G183gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(KEYINPUT26), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(G190gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT95), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n429_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G183gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n433_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n422_), .A2(new_n443_), .B1(G169gat), .B2(G176gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G169gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n424_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(G211gat), .A2(G218gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G211gat), .A2(G218gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT89), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT21), .ZN(new_n452_));
  AND2_X1   g251(.A1(G197gat), .A2(G204gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G197gat), .A2(G204gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G197gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n272_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G197gat), .A2(G204gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(KEYINPUT21), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n461_));
  INV_X1    g260(.A(new_n450_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G211gat), .A2(G218gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n453_), .A2(new_n454_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT21), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n419_), .B1(new_n448_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT25), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n469_), .A2(KEYINPUT77), .A3(KEYINPUT78), .A4(G183gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n442_), .A2(KEYINPUT25), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(G183gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT77), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT78), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n471_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n432_), .A2(new_n434_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n429_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n467_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n460_), .A2(new_n466_), .A3(KEYINPUT90), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT22), .ZN(new_n485_));
  OAI21_X1  g284(.A(G169gat), .B1(new_n485_), .B2(KEYINPUT79), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(new_n423_), .A3(KEYINPUT22), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .A4(new_n424_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n488_), .A3(new_n424_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT80), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n444_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .A4(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n418_), .B1(new_n468_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n483_), .A2(new_n484_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n477_), .B1(new_n476_), .B2(new_n436_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n480_), .B1(new_n498_), .B2(new_n470_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n493_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n419_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n429_), .A2(new_n440_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n467_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n417_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n415_), .B1(new_n496_), .B2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n444_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n476_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n476_), .B1(new_n469_), .B2(G183gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT78), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n470_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n500_), .B1(new_n513_), .B2(new_n479_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n460_), .A2(new_n466_), .A3(KEYINPUT90), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT90), .B1(new_n460_), .B2(new_n466_), .ZN(new_n516_));
  OAI22_X1  g315(.A1(new_n508_), .A2(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n517_), .A2(new_n505_), .A3(KEYINPUT20), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n518_), .A2(new_n495_), .A3(new_n414_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n409_), .B1(new_n507_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n467_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n460_), .A2(new_n466_), .A3(KEYINPUT92), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n394_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n521_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G78gat), .B(G106gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT93), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n497_), .A2(new_n521_), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n531_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n497_), .A2(new_n521_), .A3(new_n532_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n528_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n537_), .A3(KEYINPUT94), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n540_), .B1(new_n394_), .B2(KEYINPUT29), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G22gat), .B(G50gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n543_));
  INV_X1    g342(.A(new_n540_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n380_), .A2(new_n543_), .A3(new_n385_), .A4(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n542_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n539_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n541_), .A2(new_n545_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n542_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT88), .A3(new_n546_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n529_), .A2(new_n533_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT94), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n535_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n538_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n448_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n503_), .A2(KEYINPUT99), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n460_), .A2(new_n466_), .A3(KEYINPUT92), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT92), .B1(new_n460_), .B2(new_n466_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n418_), .B1(new_n565_), .B2(new_n502_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n468_), .A2(new_n494_), .A3(new_n418_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n414_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n496_), .A2(new_n415_), .A3(new_n506_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT27), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n555_), .A2(new_n530_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n572_), .A2(new_n534_), .A3(new_n546_), .A4(new_n552_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n520_), .A2(new_n558_), .A3(new_n571_), .A4(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G15gat), .B(G43gat), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n508_), .B2(new_n514_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n481_), .A2(KEYINPUT30), .A3(new_n493_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G227gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT81), .Z(new_n581_));
  XNOR2_X1  g380(.A(G71gat), .B(G99gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n576_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n508_), .A2(new_n514_), .A3(new_n577_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT30), .B1(new_n481_), .B2(new_n493_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n583_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n575_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n587_), .A2(new_n592_), .A3(KEYINPUT82), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT83), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT83), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n587_), .A2(new_n592_), .A3(KEYINPUT82), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n360_), .B(KEYINPUT31), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n587_), .A2(new_n592_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT82), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n604_));
  AOI211_X1 g403(.A(new_n408_), .B(new_n574_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n414_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n518_), .A2(new_n495_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n565_), .A2(new_n502_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n417_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n567_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n608_), .B1(new_n611_), .B2(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n408_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n380_), .A2(new_n385_), .A3(new_n360_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n614_), .A2(new_n386_), .A3(new_n399_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n400_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT4), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n388_), .A2(new_n389_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n406_), .B2(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n401_), .A2(new_n390_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n346_), .B1(new_n624_), .B2(KEYINPUT33), .ZN(new_n625_));
  INV_X1    g424(.A(new_n391_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n617_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n627_), .A2(KEYINPUT33), .A3(new_n346_), .A4(new_n405_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n414_), .B1(new_n518_), .B2(new_n495_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n628_), .A2(new_n570_), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n613_), .B1(new_n625_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n558_), .A2(new_n573_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n520_), .A2(new_n571_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n408_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n634_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT84), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n601_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n599_), .A2(new_n600_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n598_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n594_), .A2(new_n596_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n603_), .A2(KEYINPUT84), .A3(new_n604_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n605_), .B1(new_n641_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n341_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT34), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT35), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n248_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n658_));
  OAI22_X1  g457(.A1(new_n321_), .A2(new_n248_), .B1(KEYINPUT35), .B2(new_n653_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n248_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n656_), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n293_), .A2(new_n657_), .B1(new_n655_), .B2(new_n654_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(KEYINPUT36), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n664_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n667_), .B(KEYINPUT36), .Z(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT37), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n670_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n660_), .A2(new_n664_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n671_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT37), .B1(new_n677_), .B2(new_n669_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(G231gat), .A2(G233gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n308_), .B(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n254_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n320_), .A2(new_n680_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n308_), .B1(G231gat), .B2(G233gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n253_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(G127gat), .B(G155gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT16), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(G183gat), .ZN(new_n689_));
  INV_X1    g488(.A(G211gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT17), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT74), .B1(new_n686_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n686_), .A2(new_n692_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT17), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n691_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(new_n686_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n693_), .B1(new_n697_), .B2(KEYINPUT74), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n679_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n651_), .A2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n700_), .A2(G1gat), .A3(new_n639_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n701_), .A2(KEYINPUT38), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(KEYINPUT38), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n670_), .A2(new_n673_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n650_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n698_), .A3(new_n340_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G1gat), .B1(new_n706_), .B2(new_n639_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n702_), .A2(new_n703_), .A3(new_n707_), .ZN(G1324gat));
  OAI21_X1  g507(.A(G8gat), .B1(new_n706_), .B2(new_n638_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT39), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n637_), .A2(new_n295_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n700_), .B2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n706_), .B2(new_n649_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT41), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n700_), .A2(G15gat), .A3(new_n649_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1326gat));
  NOR2_X1   g516(.A1(new_n706_), .A2(new_n635_), .ZN(new_n718_));
  INV_X1    g517(.A(G22gat), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n718_), .A2(KEYINPUT100), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT100), .B1(new_n718_), .B2(new_n719_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(KEYINPUT42), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT42), .B1(new_n720_), .B2(new_n721_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n634_), .A2(new_n719_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n722_), .A2(new_n723_), .B1(new_n700_), .B2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT101), .Z(G1327gat));
  INV_X1    g525(.A(new_n704_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n698_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n651_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G29gat), .B1(new_n730_), .B2(new_n408_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n732_));
  INV_X1    g531(.A(new_n679_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n648_), .A2(new_n647_), .B1(new_n636_), .B2(new_n640_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n732_), .B(new_n733_), .C1(new_n734_), .C2(new_n605_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT102), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n649_), .A2(new_n641_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n605_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n732_), .A4(new_n733_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n650_), .B2(new_n679_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n341_), .A2(new_n698_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(KEYINPUT44), .A3(new_n744_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n408_), .A2(G29gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n731_), .B1(new_n749_), .B2(new_n750_), .ZN(G1328gat));
  OR2_X1    g550(.A1(new_n638_), .A2(KEYINPUT105), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n638_), .A2(KEYINPUT105), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(G36gat), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n729_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT107), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n637_), .A3(new_n748_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT103), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n747_), .A2(new_n764_), .A3(new_n637_), .A4(new_n748_), .ZN(new_n765_));
  AND4_X1   g564(.A1(KEYINPUT104), .A2(new_n763_), .A3(G36gat), .A4(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(G36gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n762_), .B2(KEYINPUT103), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT104), .B1(new_n768_), .B2(new_n765_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT46), .B(new_n761_), .C1(new_n766_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1329gat));
  NOR3_X1   g573(.A1(new_n729_), .A2(G43gat), .A3(new_n649_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n603_), .A2(new_n604_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n749_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(G43gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g578(.A1(new_n730_), .A2(new_n315_), .A3(new_n634_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n749_), .A2(new_n634_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n315_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT108), .ZN(G1331gat));
  INV_X1    g582(.A(new_n339_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n281_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n705_), .A2(new_n698_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT110), .B1(new_n408_), .B2(G57gat), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G57gat), .B1(new_n788_), .B2(KEYINPUT110), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n739_), .A2(new_n785_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n679_), .A2(new_n698_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT109), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n788_), .A2(new_n408_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n789_), .B1(new_n794_), .B2(new_n795_), .ZN(G1332gat));
  OAI21_X1  g595(.A(G64gat), .B1(new_n786_), .B2(new_n755_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT48), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n755_), .A2(G64gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n794_), .B2(new_n799_), .ZN(G1333gat));
  OAI21_X1  g599(.A(G71gat), .B1(new_n786_), .B2(new_n649_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT49), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n649_), .A2(G71gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n794_), .B2(new_n803_), .ZN(G1334gat));
  OAI21_X1  g603(.A(G78gat), .B1(new_n786_), .B2(new_n635_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT50), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n635_), .A2(G78gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n794_), .B2(new_n807_), .ZN(G1335gat));
  NOR3_X1   g607(.A1(new_n698_), .A2(new_n281_), .A3(new_n784_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n743_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810_), .B2(new_n639_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n790_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n728_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n813_), .A2(G85gat), .A3(new_n639_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT111), .Z(G1336gat));
  AND4_X1   g615(.A1(new_n214_), .A2(new_n743_), .A3(new_n754_), .A4(new_n809_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n813_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G92gat), .B1(new_n818_), .B2(new_n637_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1337gat));
  OAI21_X1  g619(.A(G99gat), .B1(new_n810_), .B2(new_n649_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n208_), .A3(new_n776_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g623(.A(G106gat), .B1(new_n810_), .B2(new_n635_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT52), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n818_), .A2(new_n209_), .A3(new_n634_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n329_), .A2(new_n338_), .A3(new_n278_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n266_), .A2(new_n256_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n248_), .A2(new_n254_), .B1(KEYINPUT70), .B2(KEYINPUT12), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n263_), .A2(KEYINPUT112), .A3(new_n256_), .A4(new_n266_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n259_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n267_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n833_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(new_n264_), .A3(new_n263_), .A4(new_n840_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n837_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT114), .B1(new_n846_), .B2(new_n276_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n831_), .B1(new_n847_), .B2(KEYINPUT56), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n833_), .A2(new_n834_), .A3(new_n259_), .A4(new_n841_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n842_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n844_), .A2(new_n264_), .A3(new_n263_), .A4(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n841_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n275_), .B1(new_n853_), .B2(new_n837_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n849_), .B1(new_n854_), .B2(KEYINPUT114), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n330_), .A2(new_n310_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n336_), .A2(new_n309_), .A3(new_n331_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n328_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n327_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n860_), .A2(new_n862_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n704_), .B1(new_n856_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n278_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n846_), .A2(new_n276_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n849_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n276_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n679_), .B1(new_n870_), .B2(KEYINPUT58), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872_));
  INV_X1    g671(.A(new_n869_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n276_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n875_), .B2(new_n866_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n865_), .A2(KEYINPUT57), .B1(new_n871_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n863_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n704_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT115), .B(new_n878_), .C1(new_n879_), .C2(new_n704_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n877_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n698_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n699_), .A2(new_n887_), .A3(new_n281_), .A4(new_n339_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n281_), .A2(new_n339_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n791_), .B2(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n886_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n886_), .A2(KEYINPUT116), .A3(new_n892_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n574_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n776_), .A2(new_n408_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n896_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n877_), .A2(new_n880_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT118), .B1(new_n901_), .B2(new_n885_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n891_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(KEYINPUT118), .A3(new_n885_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n898_), .A2(KEYINPUT59), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n900_), .A2(KEYINPUT59), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n355_), .B1(new_n907_), .B2(new_n784_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT116), .B1(new_n886_), .B2(new_n892_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n894_), .B(new_n891_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(KEYINPUT117), .A3(new_n899_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n339_), .A2(G113gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n910_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n830_), .B1(new_n908_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n900_), .A2(KEYINPUT59), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n905_), .A2(new_n906_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n919_), .A2(new_n784_), .A3(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT119), .B(new_n916_), .C1(new_n921_), .C2(new_n355_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n922_), .ZN(G1340gat));
  AOI21_X1  g722(.A(new_n353_), .B1(new_n907_), .B2(new_n282_), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT60), .B1(new_n282_), .B2(new_n353_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(KEYINPUT60), .B2(new_n353_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n910_), .A2(new_n914_), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT120), .B1(new_n924_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n919_), .A2(new_n282_), .A3(new_n920_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n930_), .B(new_n927_), .C1(new_n931_), .C2(new_n353_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(G1341gat));
  AND3_X1   g732(.A1(new_n907_), .A2(G127gat), .A3(new_n698_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n910_), .A2(new_n914_), .A3(new_n698_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n350_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n935_), .A2(KEYINPUT121), .A3(new_n350_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n934_), .B1(new_n938_), .B2(new_n939_), .ZN(G1342gat));
  AND2_X1   g739(.A1(new_n907_), .A2(new_n733_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n910_), .A2(new_n914_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n704_), .A2(new_n348_), .ZN(new_n943_));
  OAI22_X1  g742(.A1(new_n941_), .A2(new_n348_), .B1(new_n942_), .B2(new_n943_), .ZN(G1343gat));
  AND2_X1   g743(.A1(new_n913_), .A2(new_n649_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n754_), .A2(new_n639_), .A3(new_n635_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(new_n374_), .A3(new_n784_), .ZN(new_n949_));
  OAI21_X1  g748(.A(G141gat), .B1(new_n947_), .B2(new_n339_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1344gat));
  XNOR2_X1  g750(.A(KEYINPUT122), .B(G148gat), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n953_), .B1(new_n948_), .B2(new_n282_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n947_), .A2(new_n281_), .A3(new_n952_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(new_n955_), .ZN(G1345gat));
  XNOR2_X1  g755(.A(KEYINPUT61), .B(G155gat), .ZN(new_n957_));
  OR3_X1    g756(.A1(new_n947_), .A2(new_n885_), .A3(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n947_), .B2(new_n885_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1346gat));
  OAI21_X1  g759(.A(G162gat), .B1(new_n947_), .B2(new_n679_), .ZN(new_n961_));
  OR2_X1    g760(.A1(new_n727_), .A2(G162gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n947_), .B2(new_n962_), .ZN(G1347gat));
  AOI21_X1  g762(.A(new_n634_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n755_), .A2(new_n408_), .A3(new_n649_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(G169gat), .B1(new_n966_), .B2(new_n339_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n968_));
  OR2_X1    g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n964_), .A2(new_n445_), .A3(new_n784_), .A4(new_n965_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n967_), .A2(new_n968_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n969_), .A2(new_n970_), .A3(new_n971_), .ZN(G1348gat));
  OAI21_X1  g771(.A(new_n424_), .B1(new_n966_), .B2(new_n281_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n911_), .A2(new_n912_), .A3(new_n634_), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n974_), .A2(G176gat), .A3(new_n282_), .A4(new_n965_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n976_), .B(new_n977_), .ZN(G1349gat));
  AND2_X1   g777(.A1(new_n965_), .A2(new_n698_), .ZN(new_n979_));
  AND3_X1   g778(.A1(new_n964_), .A2(new_n474_), .A3(new_n979_), .ZN(new_n980_));
  AOI21_X1  g779(.A(KEYINPUT124), .B1(new_n974_), .B2(new_n979_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n981_), .A2(G183gat), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n974_), .A2(KEYINPUT124), .A3(new_n979_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n980_), .B1(new_n982_), .B2(new_n983_), .ZN(G1350gat));
  OAI21_X1  g783(.A(G190gat), .B1(new_n966_), .B2(new_n679_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n704_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n985_), .B1(new_n966_), .B2(new_n986_), .ZN(G1351gat));
  NOR3_X1   g786(.A1(new_n755_), .A2(new_n408_), .A3(new_n635_), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n913_), .A2(new_n649_), .A3(new_n988_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n989_), .A2(new_n339_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(new_n456_), .ZN(G1352gat));
  NOR2_X1   g790(.A1(new_n989_), .A2(new_n281_), .ZN(new_n992_));
  NOR2_X1   g791(.A1(new_n272_), .A2(KEYINPUT125), .ZN(new_n993_));
  XOR2_X1   g792(.A(new_n992_), .B(new_n993_), .Z(G1353gat));
  AND2_X1   g793(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n995_));
  NOR2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  NOR4_X1   g795(.A1(new_n989_), .A2(new_n885_), .A3(new_n995_), .A4(new_n996_), .ZN(new_n997_));
  OAI21_X1  g796(.A(new_n996_), .B1(new_n989_), .B2(new_n885_), .ZN(new_n998_));
  OR2_X1    g797(.A1(new_n998_), .A2(KEYINPUT126), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n998_), .A2(KEYINPUT126), .ZN(new_n1000_));
  AOI21_X1  g799(.A(new_n997_), .B1(new_n999_), .B2(new_n1000_), .ZN(G1354gat));
  OAI21_X1  g800(.A(G218gat), .B1(new_n989_), .B2(new_n679_), .ZN(new_n1002_));
  OR2_X1    g801(.A1(new_n727_), .A2(G218gat), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1002_), .B1(new_n989_), .B2(new_n1003_), .ZN(G1355gat));
endmodule


