//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT82), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT3), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT3), .B1(new_n205_), .B2(new_n206_), .ZN(new_n208_));
  OAI22_X1  g007(.A1(new_n207_), .A2(new_n208_), .B1(KEYINPUT83), .B2(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n203_), .B(new_n204_), .C1(new_n209_), .C2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(new_n206_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n202_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n204_), .B(KEYINPUT1), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n214_), .B(new_n210_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT79), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n220_), .A2(new_n221_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT80), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n220_), .A2(new_n221_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n213_), .B(new_n218_), .C1(new_n227_), .C2(new_n224_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n226_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT99), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n226_), .B2(KEYINPUT4), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT100), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n226_), .A2(new_n228_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT101), .B1(new_n238_), .B2(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(KEYINPUT101), .A3(new_n236_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G57gat), .B(G85gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(G1gat), .B(G29gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n236_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n230_), .B(new_n232_), .C1(KEYINPUT4), .C2(new_n226_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n229_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n239_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n241_), .B(new_n249_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT97), .ZN(new_n256_));
  OR2_X1    g055(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT24), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n259_), .A2(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT24), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(G183gat), .B2(G190gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(G183gat), .A3(G190gat), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT78), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT78), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT22), .B(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(G176gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n264_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT96), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n279_), .A3(new_n264_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n269_), .A2(KEYINPUT76), .ZN(new_n281_));
  INV_X1    g080(.A(new_n268_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n269_), .A2(KEYINPUT76), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n278_), .B(new_n280_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n273_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G204gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT88), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT88), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G204gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n292_), .A3(G197gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n289_), .B2(G197gat), .ZN(new_n295_));
  INV_X1    g094(.A(G197gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G211gat), .B(G218gat), .Z(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(KEYINPUT21), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302_));
  AND4_X1   g101(.A1(new_n302_), .A2(new_n293_), .A3(new_n295_), .A4(new_n297_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT89), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT88), .B(G204gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(G197gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n290_), .A2(new_n292_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(KEYINPUT89), .A3(new_n296_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n289_), .A2(G197gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n303_), .B1(new_n310_), .B2(KEYINPUT21), .ZN(new_n311_));
  INV_X1    g110(.A(new_n299_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n301_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n256_), .B1(new_n288_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT20), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n264_), .B1(new_n272_), .B2(new_n286_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n276_), .B(KEYINPUT77), .ZN(new_n317_));
  OAI22_X1  g116(.A1(new_n316_), .A2(new_n317_), .B1(new_n285_), .B2(new_n266_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n315_), .B1(new_n319_), .B2(new_n313_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(KEYINPUT21), .ZN(new_n321_));
  INV_X1    g120(.A(new_n303_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n312_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n300_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n273_), .A2(new_n287_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT97), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n314_), .A2(new_n320_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G8gat), .B(G36gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G92gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT18), .B(G64gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n329_), .B1(new_n288_), .B2(new_n313_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT98), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n319_), .B2(new_n313_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n324_), .A2(KEYINPUT98), .A3(new_n318_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT20), .A4(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n327_), .A2(new_n329_), .ZN(new_n342_));
  AOI211_X1 g141(.A(KEYINPUT92), .B(new_n301_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n323_), .B2(new_n300_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n288_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n346_), .A2(KEYINPUT20), .A3(new_n338_), .A4(new_n339_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n342_), .B1(new_n329_), .B2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(KEYINPUT27), .B(new_n341_), .C1(new_n348_), .C2(new_n335_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT106), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT27), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n329_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n329_), .B2(new_n327_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n353_), .B2(new_n334_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT106), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n341_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n341_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n335_), .B1(new_n330_), .B2(new_n340_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n351_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT86), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n343_), .A2(new_n345_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n364_), .B(KEYINPUT87), .Z(new_n368_));
  NAND3_X1  g167(.A1(new_n324_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT91), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT91), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n324_), .A2(new_n371_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n362_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT93), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n324_), .A2(KEYINPUT92), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n313_), .A2(new_n344_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n366_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n364_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(new_n361_), .A3(new_n370_), .A4(new_n372_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n219_), .A2(KEYINPUT85), .A3(KEYINPUT29), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT85), .B1(new_n219_), .B2(KEYINPUT29), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G22gat), .B(G50gat), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n384_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(new_n391_), .A3(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n367_), .A2(new_n373_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT93), .A3(new_n361_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n382_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT94), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT95), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n374_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n381_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n395_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n400_), .A3(new_n361_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n382_), .A2(new_n406_), .A3(new_n397_), .A4(new_n395_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n399_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n225_), .A2(new_n223_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(new_n318_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G71gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT30), .B(G99gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n412_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n408_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n399_), .A2(new_n405_), .A3(new_n407_), .A4(new_n421_), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n255_), .B(new_n360_), .C1(new_n420_), .C2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n254_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n240_), .A2(KEYINPUT33), .A3(new_n249_), .A4(new_n241_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT104), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n234_), .A2(new_n250_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n238_), .B(KEYINPUT103), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n429_), .B(new_n247_), .C1(new_n250_), .C2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n357_), .A2(new_n358_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n428_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n432_), .A2(new_n431_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT104), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n330_), .A2(new_n340_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT105), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT105), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n353_), .B2(new_n437_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n255_), .B(new_n439_), .C1(new_n438_), .C2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n408_), .A2(new_n421_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n423_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447_));
  XOR2_X1   g246(.A(G183gat), .B(G211gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(G127gat), .B(G155gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n447_), .B1(new_n452_), .B2(KEYINPUT17), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454_));
  INV_X1    g253(.A(G1gat), .ZN(new_n455_));
  INV_X1    g254(.A(G8gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT14), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G8gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n453_), .B(new_n460_), .Z(new_n461_));
  NAND2_X1  g260(.A1(G231gat), .A2(G233gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(G57gat), .A2(G64gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT11), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G57gat), .A2(G64gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470_));
  INV_X1    g269(.A(G78gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G71gat), .ZN(new_n472_));
  INV_X1    g271(.A(G71gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G78gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G57gat), .A2(G64gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G57gat), .A2(G64gat), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT66), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n478_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n465_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n452_), .A2(KEYINPUT17), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n480_), .A2(new_n487_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n463_), .A2(new_n490_), .A3(new_n464_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT71), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT35), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500_));
  OR2_X1    g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT9), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT10), .B(G99gat), .Z(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n504_), .A2(new_n507_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT8), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT65), .B1(new_n508_), .B2(new_n509_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT6), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  NAND3_X1  g321(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(new_n518_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n513_), .B1(new_n525_), .B2(new_n503_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT64), .B(KEYINPUT8), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n502_), .A3(new_n501_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n512_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G43gat), .B(G50gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G29gat), .B(G36gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n512_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n525_), .A2(new_n503_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT8), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  INV_X1    g337(.A(new_n529_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT68), .B1(new_n526_), .B2(new_n529_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n535_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n533_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n500_), .B(new_n534_), .C1(new_n542_), .C2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n498_), .A2(KEYINPUT35), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n499_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n526_), .A2(KEYINPUT68), .A3(new_n529_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n512_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT72), .B1(new_n551_), .B2(new_n544_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n552_), .A2(KEYINPUT35), .A3(new_n498_), .A4(new_n534_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT36), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n548_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT36), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n494_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT74), .B(new_n494_), .C1(new_n559_), .C2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n548_), .A2(new_n553_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n561_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n548_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(KEYINPUT37), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT73), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n570_), .A2(new_n574_), .A3(KEYINPUT37), .A4(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n446_), .A2(new_n493_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n447_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n479_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n485_), .A2(new_n478_), .A3(new_n486_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT67), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(G230gat), .ZN(new_n585_));
  INV_X1    g384(.A(G233gat), .ZN(new_n586_));
  OAI22_X1  g385(.A1(new_n584_), .A2(new_n530_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n490_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n583_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT67), .B1(new_n581_), .B2(new_n582_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n530_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n585_), .A2(new_n586_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n530_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n537_), .A2(new_n539_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n583_), .A2(new_n580_), .B1(new_n598_), .B2(new_n512_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G176gat), .B(G204gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n601_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT13), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n460_), .A2(new_n533_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n544_), .B2(new_n460_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n460_), .A2(new_n533_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n616_), .B2(new_n611_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n614_), .A2(new_n617_), .A3(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n610_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n579_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n455_), .A3(new_n255_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  INV_X1    g428(.A(new_n626_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n559_), .A2(new_n563_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT107), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n446_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n420_), .A2(new_n422_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n255_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n360_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n443_), .A2(new_n444_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n633_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT108), .A3(new_n641_), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n493_), .B(new_n630_), .C1(new_n634_), .C2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(new_n255_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n629_), .B1(new_n455_), .B2(new_n644_), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n634_), .A2(new_n642_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n492_), .A3(new_n626_), .A4(new_n360_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G8gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT109), .B(KEYINPUT39), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n627_), .A2(new_n456_), .A3(new_n360_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(G8gat), .A3(new_n649_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n651_), .A2(KEYINPUT40), .A3(new_n652_), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  INV_X1    g457(.A(G15gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n627_), .A2(new_n659_), .A3(new_n421_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n643_), .A2(new_n421_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n661_), .B2(G15gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n627_), .A2(new_n665_), .A3(new_n408_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n643_), .A2(new_n408_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(G22gat), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT42), .B(new_n665_), .C1(new_n643_), .C2(new_n408_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1327gat));
  INV_X1    g470(.A(KEYINPUT111), .ZN(new_n672_));
  INV_X1    g471(.A(new_n632_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n493_), .B(new_n673_), .C1(new_n423_), .C2(new_n445_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n674_), .B2(new_n630_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n492_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n676_), .A2(KEYINPUT111), .A3(new_n626_), .A4(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n255_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n577_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n681_), .B1(new_n640_), .B2(new_n684_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT43), .B(new_n577_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n493_), .B(new_n626_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n640_), .A2(new_n681_), .A3(new_n578_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n683_), .B1(new_n639_), .B2(new_n638_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n681_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n493_), .A4(new_n626_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n689_), .A2(new_n255_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n680_), .B1(new_n694_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n689_), .A2(new_n360_), .A3(new_n693_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n675_), .A2(new_n698_), .A3(new_n360_), .A4(new_n677_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT45), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n700_), .A3(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND4_X1  g504(.A1(new_n689_), .A2(new_n693_), .A3(G43gat), .A4(new_n421_), .ZN(new_n706_));
  INV_X1    g505(.A(G43gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n678_), .B2(new_n419_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g509(.A1(G50gat), .A2(new_n689_), .A3(new_n408_), .A4(new_n693_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G50gat), .B1(new_n679_), .B2(new_n408_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n625_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n609_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n579_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n255_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n646_), .A2(new_n492_), .A3(new_n715_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n255_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g519(.A(G64gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n721_), .A3(new_n360_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n360_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G64gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT48), .B(new_n721_), .C1(new_n718_), .C2(new_n360_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n473_), .A3(new_n421_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n718_), .A2(new_n421_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G71gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT49), .B(new_n473_), .C1(new_n718_), .C2(new_n421_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1334gat));
  AND2_X1   g532(.A1(new_n715_), .A2(new_n408_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n579_), .A2(new_n471_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n718_), .A2(new_n408_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G78gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT50), .B(new_n471_), .C1(new_n718_), .C2(new_n408_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n674_), .A2(new_n714_), .A3(new_n609_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n255_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n692_), .A2(KEYINPUT112), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n690_), .B(new_n744_), .C1(new_n691_), .C2(new_n681_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n743_), .A2(new_n493_), .A3(new_n745_), .A4(new_n715_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n636_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n747_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g547(.A(G92gat), .B1(new_n741_), .B2(new_n360_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n746_), .A2(new_n637_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n746_), .B2(new_n419_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n505_), .A3(new_n421_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n756_), .A3(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1338gat));
  NAND3_X1  g557(.A1(new_n741_), .A2(new_n506_), .A3(new_n408_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n692_), .A2(new_n493_), .A3(new_n734_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G106gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G106gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n759_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n360_), .A2(new_n422_), .A3(new_n636_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n595_), .A2(new_n600_), .A3(new_n607_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n612_), .A2(new_n615_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n613_), .B1(new_n616_), .B2(new_n611_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n621_), .A3(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(new_n624_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n773_), .A2(new_n777_), .A3(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n490_), .A2(KEYINPUT12), .ZN(new_n783_));
  OAI22_X1  g582(.A1(new_n599_), .A2(KEYINPUT12), .B1(new_n542_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n596_), .B1(new_n784_), .B2(new_n597_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n784_), .B2(new_n587_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT55), .A4(new_n594_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n606_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n606_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT56), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n782_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT58), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n782_), .A2(new_n796_), .A3(new_n793_), .A4(new_n791_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n577_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n625_), .B1(new_n601_), .B2(new_n607_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n789_), .B2(new_n606_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(KEYINPUT56), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n801_), .B(new_n790_), .C1(new_n789_), .C2(new_n606_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n792_), .A2(KEYINPUT113), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n790_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n792_), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n807_), .A2(KEYINPUT114), .A3(new_n800_), .A4(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n608_), .A2(new_n777_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n805_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n632_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n798_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n492_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n609_), .A2(new_n577_), .A3(new_n492_), .A4(new_n625_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n817_), .B(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n771_), .B(new_n772_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT117), .B(new_n772_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n770_), .A2(new_n820_), .B1(new_n821_), .B2(KEYINPUT59), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n820_), .A2(new_n770_), .A3(KEYINPUT59), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n625_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n822_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n816_), .A2(new_n819_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n772_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n829_), .B2(new_n625_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n769_), .B1(new_n827_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n770_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n835_), .B(new_n825_), .C1(new_n836_), .C2(new_n834_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT119), .A3(new_n830_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(new_n829_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n609_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n840_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n822_), .A2(new_n823_), .A3(new_n609_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n840_), .B2(new_n492_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n822_), .A2(new_n823_), .A3(new_n493_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n822_), .A2(new_n823_), .A3(new_n849_), .A4(new_n577_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n829_), .B2(new_n641_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(G1343gat));
  INV_X1    g653(.A(new_n420_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n360_), .A2(new_n636_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n828_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n625_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n205_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n609_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n206_), .ZN(G1345gat));
  AND2_X1   g660(.A1(new_n828_), .A2(new_n855_), .ZN(new_n862_));
  INV_X1    g661(.A(G155gat), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n492_), .A4(new_n856_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G155gat), .B1(new_n857_), .B2(new_n493_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1346gat));
  NAND4_X1  g668(.A1(new_n862_), .A2(G162gat), .A3(new_n684_), .A4(new_n856_), .ZN(new_n870_));
  INV_X1    g669(.A(G162gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n857_), .B2(new_n641_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(KEYINPUT122), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1347gat));
  NOR3_X1   g676(.A1(new_n637_), .A2(new_n255_), .A3(new_n422_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n828_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n714_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n714_), .A2(new_n274_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT123), .ZN(new_n886_));
  OAI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n879_), .B2(new_n886_), .ZN(G1348gat));
  NOR2_X1   g686(.A1(new_n879_), .A2(new_n609_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT124), .B(G176gat), .Z(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1349gat));
  NAND2_X1  g689(.A1(new_n880_), .A2(new_n492_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n258_), .B1(new_n257_), .B2(KEYINPUT125), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT125), .A2(G183gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n891_), .B2(new_n894_), .ZN(G1350gat));
  NAND3_X1  g694(.A1(new_n880_), .A2(new_n260_), .A3(new_n633_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G190gat), .B1(new_n879_), .B2(new_n577_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n637_), .A2(new_n255_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n862_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT126), .B(G197gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n714_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n900_), .B2(new_n625_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1352gat));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(G204gat), .C1(new_n900_), .C2(new_n609_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n901_), .A2(new_n610_), .A3(new_n290_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n292_), .A2(KEYINPUT127), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1353gat));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n901_), .B(new_n492_), .C1(new_n912_), .C2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n900_), .A2(new_n493_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n912_), .ZN(G1354gat));
  INV_X1    g715(.A(G218gat), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n900_), .A2(new_n917_), .A3(new_n577_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n901_), .A2(new_n633_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(new_n919_), .ZN(G1355gat));
endmodule


