//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT1), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n208_), .B(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(KEYINPUT83), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT2), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n202_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(new_n203_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n210_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n221_), .B(KEYINPUT28), .Z(new_n222_));
  XOR2_X1   g021(.A(G22gat), .B(G50gat), .Z(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G197gat), .B(G204gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(G211gat), .B(G218gat), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT21), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n225_), .A3(KEYINPUT21), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT84), .B(KEYINPUT29), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n219_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G228gat), .ZN(new_n236_));
  INV_X1    g035(.A(G233gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  OAI221_X1 g038(.A(new_n233_), .B1(new_n236_), .B2(new_n237_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n224_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n241_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n243_), .A3(new_n223_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n222_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n222_), .A3(new_n249_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G71gat), .B(G99gat), .Z(new_n253_));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G15gat), .B(G43gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT82), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n255_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT23), .ZN(new_n261_));
  OR2_X1    g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n262_), .A2(KEYINPUT24), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n266_), .A2(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT78), .B(G183gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT79), .B(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT26), .ZN(new_n276_));
  OR2_X1    g075(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n273_), .A2(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT22), .B(G169gat), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT81), .ZN(new_n283_));
  INV_X1    g082(.A(new_n275_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n271_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n261_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n265_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT30), .B1(new_n279_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(KEYINPUT30), .A3(new_n287_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n259_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n290_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n292_), .A2(new_n258_), .A3(new_n288_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT31), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n258_), .B1(new_n292_), .B2(new_n288_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n289_), .A2(new_n259_), .A3(new_n290_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n294_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n297_), .B1(new_n294_), .B2(new_n301_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n251_), .B(new_n252_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n294_), .A2(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n297_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n252_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n308_), .B(new_n302_), .C1(new_n309_), .C2(new_n250_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n231_), .A2(new_n232_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT25), .B(G183gat), .Z(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT26), .B(G190gat), .Z(new_n318_));
  OAI211_X1 g117(.A(new_n264_), .B(new_n266_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n265_), .B(KEYINPUT86), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n282_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n316_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(KEYINPUT20), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n316_), .B1(new_n279_), .B2(new_n287_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n325_), .B(KEYINPUT85), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n279_), .A2(new_n287_), .A3(new_n316_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n319_), .A2(new_n322_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n233_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n315_), .B1(new_n329_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT87), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n329_), .A2(new_n336_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n315_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n329_), .A2(new_n336_), .A3(new_n315_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT87), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n332_), .A2(new_n335_), .A3(new_n331_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n323_), .A2(KEYINPUT20), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT92), .ZN(new_n349_));
  INV_X1    g148(.A(new_n328_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n323_), .A2(new_n351_), .A3(KEYINPUT20), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n347_), .B1(new_n353_), .B2(new_n325_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n341_), .B1(new_n354_), .B2(new_n340_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT27), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n219_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n307_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n219_), .A2(new_n297_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n219_), .A2(new_n297_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT89), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  NOR4_X1   g166(.A1(new_n219_), .A2(new_n367_), .A3(KEYINPUT4), .A4(new_n297_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n361_), .B(new_n363_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n359_), .A2(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G1gat), .B(G29gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT0), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(KEYINPUT90), .Z(new_n375_));
  XNOR2_X1  g174(.A(G57gat), .B(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n357_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n311_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n303_), .A2(new_n304_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n366_), .A2(new_n368_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(KEYINPUT91), .A3(new_n362_), .A4(new_n361_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n377_), .B1(new_n370_), .B2(new_n363_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n361_), .B(new_n362_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n380_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n369_), .A2(new_n371_), .A3(KEYINPUT33), .A4(new_n377_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n392_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n344_), .B1(KEYINPUT87), .B2(new_n337_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n344_), .A2(KEYINPUT87), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n342_), .A2(KEYINPUT88), .A3(new_n345_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n340_), .A2(KEYINPUT32), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n353_), .A2(new_n325_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n403_), .B(new_n405_), .C1(new_n406_), .C2(new_n347_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n339_), .A2(new_n404_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT93), .B1(new_n354_), .B2(new_n404_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n407_), .A2(new_n381_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n385_), .B1(new_n402_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n384_), .B1(new_n411_), .B2(new_n311_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G113gat), .B(G141gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT77), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G169gat), .B(G197gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G229gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(G1gat), .ZN(new_n419_));
  INV_X1    g218(.A(G8gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G22gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G15gat), .ZN(new_n423_));
  INV_X1    g222(.A(G15gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G22gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT73), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G8gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n426_), .A2(KEYINPUT73), .ZN(new_n430_));
  INV_X1    g229(.A(new_n428_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(KEYINPUT73), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G43gat), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G29gat), .B(G36gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT68), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(KEYINPUT68), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n436_), .A2(KEYINPUT68), .ZN(new_n441_));
  INV_X1    g240(.A(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n429_), .A2(new_n444_), .A3(new_n433_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n418_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT75), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n438_), .A2(new_n439_), .A3(new_n435_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n442_), .B1(new_n441_), .B2(new_n437_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT15), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT15), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n440_), .A2(new_n454_), .A3(new_n443_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n453_), .A2(new_n455_), .A3(new_n433_), .A4(new_n429_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n418_), .B(KEYINPUT76), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n446_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n448_), .B2(KEYINPUT75), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n417_), .B1(new_n450_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n446_), .A2(new_n447_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n418_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n417_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n449_), .A3(new_n458_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n413_), .A2(KEYINPUT94), .A3(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G71gat), .B(G78gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G64gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G57gat), .ZN(new_n473_));
  INV_X1    g272(.A(G57gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G64gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT11), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n473_), .A2(new_n475_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n470_), .B1(new_n478_), .B2(KEYINPUT11), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(G85gat), .A2(G92gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT9), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT65), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n483_), .A2(new_n485_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n485_), .A2(new_n488_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n489_), .A2(new_n490_), .A3(new_n494_), .A4(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n483_), .A2(new_n488_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n501_), .B1(new_n505_), .B2(new_n494_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n500_), .B1(new_n506_), .B2(KEYINPUT8), .ZN(new_n507_));
  XOR2_X1   g306(.A(G85gat), .B(G92gat), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n497_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT66), .A3(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n509_), .B1(new_n516_), .B2(new_n494_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n482_), .B1(new_n507_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT64), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n490_), .A2(new_n494_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n525_));
  AND2_X1   g324(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n495_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n508_), .A2(new_n525_), .B1(new_n527_), .B2(new_n497_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n514_), .A2(new_n531_), .A3(new_n491_), .A4(new_n502_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n508_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n524_), .A2(new_n528_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n514_), .A2(KEYINPUT66), .A3(new_n502_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT66), .B1(new_n514_), .B2(new_n502_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n494_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n509_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n478_), .A2(new_n470_), .A3(KEYINPUT11), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n471_), .A2(new_n476_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n479_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(new_n534_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n531_), .A2(new_n491_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(new_n500_), .C1(new_n547_), .C2(new_n509_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(KEYINPUT12), .A3(new_n482_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n520_), .A2(new_n523_), .A3(new_n544_), .A4(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n482_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n543_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n522_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT5), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G176gat), .B(G204gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n561_));
  OR3_X1    g360(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT13), .B1(new_n560_), .B2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n445_), .A2(new_n540_), .A3(new_n535_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n453_), .A2(new_n548_), .A3(new_n455_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n574_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT69), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(KEYINPUT69), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n576_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n568_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n570_), .A2(new_n575_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n584_), .A2(KEYINPUT69), .A3(new_n569_), .A4(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n576_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n567_), .B(KEYINPUT36), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n582_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n582_), .A2(KEYINPUT71), .A3(new_n583_), .A4(new_n588_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n587_), .B(KEYINPUT70), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n580_), .A2(new_n581_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n568_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT72), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n591_), .A2(new_n600_), .A3(new_n592_), .A4(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT74), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n434_), .A2(new_n543_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n429_), .A2(new_n433_), .A3(new_n482_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n609_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n607_), .A2(new_n608_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n618_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n603_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624_));
  INV_X1    g423(.A(new_n468_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n412_), .B2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n469_), .A2(new_n564_), .A3(new_n623_), .A4(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n627_), .A2(G1gat), .A3(new_n382_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT38), .Z(new_n629_));
  AND2_X1   g428(.A1(new_n582_), .A2(new_n588_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n564_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(new_n625_), .A3(new_n622_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n413_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n382_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n635_), .ZN(G1324gat));
  OAI21_X1  g435(.A(G8gat), .B1(new_n634_), .B2(new_n357_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT39), .ZN(new_n638_));
  INV_X1    g437(.A(new_n357_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n420_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n638_), .B1(new_n627_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g441(.A(new_n385_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G15gat), .B1(new_n634_), .B2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT95), .B(KEYINPUT41), .Z(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n385_), .A2(new_n424_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n627_), .B2(new_n647_), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n309_), .A2(new_n250_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G22gat), .B1(new_n634_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT96), .B(KEYINPUT42), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n422_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n627_), .B2(new_n654_), .ZN(G1327gat));
  NOR2_X1   g454(.A1(new_n631_), .A2(new_n621_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n469_), .A2(new_n564_), .A3(new_n626_), .A4(new_n656_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n657_), .A2(G29gat), .A3(new_n382_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT97), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n412_), .B2(new_n602_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(KEYINPUT97), .B2(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n412_), .A2(KEYINPUT98), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n659_), .A2(KEYINPUT98), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n384_), .B(new_n664_), .C1(new_n411_), .C2(new_n311_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n602_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n632_), .A2(new_n625_), .A3(new_n621_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n382_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n667_), .A2(new_n672_), .A3(KEYINPUT44), .A4(new_n668_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n674_));
  INV_X1    g473(.A(new_n311_), .ZN(new_n675_));
  AND4_X1   g474(.A1(new_n381_), .A2(new_n407_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT88), .B1(new_n342_), .B2(new_n345_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n392_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n679_), .B2(new_n401_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n680_), .B2(new_n385_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n674_), .B1(new_n681_), .B2(new_n384_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n665_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n603_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n659_), .A2(KEYINPUT97), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n384_), .A3(new_n603_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n660_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(KEYINPUT44), .A4(new_n668_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT99), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n673_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n671_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n671_), .B2(new_n690_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n658_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n673_), .A2(new_n689_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n639_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n357_), .B(KEYINPUT101), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n697_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n657_), .A2(KEYINPUT45), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT45), .B1(new_n657_), .B2(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n696_), .B1(new_n699_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n669_), .A2(new_n670_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n690_), .A2(new_n639_), .A3(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT46), .B(new_n704_), .C1(new_n708_), .C2(new_n697_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n690_), .A2(G43gat), .A3(new_n385_), .A4(new_n707_), .ZN(new_n711_));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n657_), .B2(new_n643_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  OR3_X1    g517(.A1(new_n657_), .A2(G50gat), .A3(new_n650_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n698_), .A2(new_n720_), .A3(new_n649_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n698_), .B2(new_n649_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1331gat));
  NOR2_X1   g523(.A1(new_n564_), .A2(new_n468_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n622_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n413_), .A2(new_n631_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n413_), .A2(KEYINPUT103), .A3(new_n631_), .A4(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n382_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n413_), .A2(new_n725_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(new_n622_), .A3(new_n603_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n474_), .A3(new_n381_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1332gat));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n472_), .A3(new_n700_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n700_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G64gat), .B1(new_n732_), .B2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(KEYINPUT48), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(KEYINPUT48), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n732_), .B2(new_n643_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n735_), .A2(new_n748_), .A3(new_n385_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(new_n747_), .A3(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n735_), .A2(new_n751_), .A3(new_n649_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n730_), .A2(new_n649_), .A3(new_n731_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G78gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT105), .Z(G1335gat));
  NOR2_X1   g557(.A1(new_n726_), .A2(new_n621_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n667_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n382_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n734_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n656_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n382_), .A2(G85gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n739_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n357_), .A2(G92gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n763_), .B2(new_n767_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n760_), .B2(new_n643_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n763_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n527_), .A3(new_n385_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT106), .B(KEYINPUT51), .Z(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1338gat));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n684_), .A2(new_n687_), .A3(new_n649_), .A4(new_n759_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(KEYINPUT52), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n776_), .A2(KEYINPUT107), .A3(new_n779_), .A4(G106gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(KEYINPUT52), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n770_), .A2(new_n497_), .A3(new_n649_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT109), .B1(new_n622_), .B2(new_n468_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n621_), .A2(new_n460_), .A3(new_n790_), .A4(new_n467_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n564_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(new_n564_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n788_), .B1(new_n796_), .B2(new_n602_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n603_), .A2(new_n794_), .A3(new_n795_), .A4(KEYINPUT54), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n560_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n544_), .B1(new_n552_), .B2(KEYINPUT12), .ZN(new_n802_));
  INV_X1    g601(.A(new_n549_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n522_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n520_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT111), .A3(new_n522_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n550_), .A2(KEYINPUT55), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT12), .B1(new_n548_), .B2(new_n482_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n551_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n523_), .A4(new_n549_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n806_), .A2(new_n808_), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n558_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n809_), .A2(new_n813_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT111), .B1(new_n807_), .B2(new_n522_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n807_), .A2(KEYINPUT111), .A3(new_n522_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n557_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n801_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n466_), .B1(new_n461_), .B2(new_n457_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n446_), .A2(new_n456_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n457_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n467_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n560_), .A2(new_n561_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n630_), .B1(new_n822_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n815_), .B1(new_n814_), .B2(new_n558_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n819_), .A2(new_n818_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n550_), .B(new_n812_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT56), .B(new_n557_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n828_), .B1(new_n838_), .B2(new_n801_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT112), .B(new_n833_), .C1(new_n839_), .C2(new_n630_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n467_), .A2(new_n559_), .A3(new_n825_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(KEYINPUT113), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT58), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n845_), .A2(new_n848_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n840_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n622_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(KEYINPUT116), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(KEYINPUT116), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n800_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n639_), .A2(new_n310_), .A3(new_n382_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(KEYINPUT114), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n832_), .A2(new_n849_), .A3(new_n859_), .A4(new_n840_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n621_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n856_), .B1(new_n861_), .B2(new_n799_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n862_), .A2(new_n863_), .A3(KEYINPUT59), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n862_), .B2(KEYINPUT59), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n857_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n625_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n625_), .A2(G113gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n862_), .B2(new_n868_), .ZN(G1340gat));
  OAI21_X1  g668(.A(G120gat), .B1(new_n866_), .B2(new_n564_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n862_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n872_));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n632_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n870_), .A2(new_n876_), .ZN(G1341gat));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n866_), .A2(new_n878_), .A3(new_n622_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n862_), .B2(new_n622_), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT117), .Z(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1342gat));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n602_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n857_), .B(new_n884_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n862_), .B2(new_n631_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(KEYINPUT118), .A3(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n858_), .A2(new_n860_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n622_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n800_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n305_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n700_), .A2(new_n382_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT119), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n894_), .A2(new_n899_), .A3(new_n895_), .A4(new_n896_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n625_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT120), .B(G141gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1344gat));
  AOI21_X1  g702(.A(new_n564_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT121), .B(G148gat), .Z(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n904_), .B(new_n906_), .ZN(G1345gat));
  AOI21_X1  g706(.A(new_n622_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT61), .B(G155gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  NAND2_X1  g709(.A1(new_n898_), .A2(new_n900_), .ZN(new_n911_));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n630_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n602_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n912_), .ZN(G1347gat));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n700_), .A2(new_n382_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n385_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n649_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n854_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n280_), .A3(new_n468_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n854_), .A2(new_n468_), .A3(new_n920_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT62), .B1(new_n923_), .B2(G169gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n916_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n926_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n928_), .A2(KEYINPUT122), .A3(new_n924_), .A4(new_n922_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1348gat));
  NAND2_X1  g729(.A1(new_n854_), .A2(new_n920_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n281_), .B1(new_n931_), .B2(new_n564_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n919_), .A2(new_n281_), .A3(new_n564_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n894_), .A2(new_n650_), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT123), .ZN(G1349gat));
  AND2_X1   g735(.A1(new_n621_), .A2(new_n317_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n919_), .A2(new_n622_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n894_), .A2(new_n650_), .A3(new_n938_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n921_), .A2(new_n937_), .B1(new_n939_), .B2(new_n271_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n931_), .B2(new_n602_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n631_), .A2(new_n318_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n931_), .B2(new_n942_), .ZN(G1351gat));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944_));
  INV_X1    g743(.A(G197gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n894_), .A2(new_n895_), .A3(new_n918_), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n944_), .B(new_n945_), .C1(new_n946_), .C2(new_n625_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n946_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n468_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n947_), .B1(new_n949_), .B2(new_n945_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n944_), .B1(new_n949_), .B2(new_n945_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1352gat));
  NAND2_X1  g751(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n948_), .A2(new_n632_), .A3(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955_));
  AOI21_X1  g754(.A(KEYINPUT126), .B1(new_n955_), .B2(G204gat), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n954_), .B(new_n956_), .Z(G1353gat));
  NOR2_X1   g756(.A1(new_n946_), .A2(new_n622_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  AND2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n958_), .B2(new_n959_), .ZN(G1354gat));
  AND3_X1   g761(.A1(new_n948_), .A2(G218gat), .A3(new_n603_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n946_), .A2(new_n631_), .ZN(new_n964_));
  OR2_X1    g763(.A1(new_n964_), .A2(KEYINPUT127), .ZN(new_n965_));
  AOI21_X1  g764(.A(G218gat), .B1(new_n964_), .B2(KEYINPUT127), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n963_), .B1(new_n965_), .B2(new_n966_), .ZN(G1355gat));
endmodule


