//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(G218gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G211gat), .ZN(new_n204_));
  INV_X1    g003(.A(G211gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G218gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT88), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT21), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT85), .B1(new_n213_), .B2(G197gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  INV_X1    g014(.A(G197gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(G204gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(G197gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n217_), .A3(KEYINPUT89), .A4(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n229_), .A2(new_n214_), .A3(new_n218_), .A4(new_n217_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n216_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n213_), .B2(G197gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n216_), .A2(G204gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT21), .B(new_n231_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  AND4_X1   g034(.A1(KEYINPUT87), .A2(new_n230_), .A3(new_n235_), .A4(new_n210_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n213_), .A2(G197gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n225_), .B1(new_n237_), .B2(KEYINPUT84), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n216_), .A2(G204gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n218_), .A3(new_n232_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n207_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT87), .B1(new_n241_), .B2(new_n230_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n224_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT90), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n246_), .A2(new_n247_), .A3(new_n254_), .A4(new_n248_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n250_), .A2(new_n253_), .A3(new_n255_), .A4(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260_));
  INV_X1    g059(.A(G169gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n257_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n246_), .A2(new_n248_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n262_), .A2(KEYINPUT24), .A3(new_n251_), .A4(new_n263_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n266_), .A2(new_n269_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n259_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n243_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n261_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n275_));
  AND2_X1   g074(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n275_), .B(new_n257_), .C1(new_n261_), .C2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n253_), .A2(new_n277_), .A3(new_n249_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n266_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n264_), .A2(new_n265_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n253_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT87), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n235_), .A2(new_n210_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n219_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n284_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n241_), .A2(KEYINPUT87), .A3(new_n230_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n283_), .A2(new_n290_), .A3(new_n224_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n274_), .A2(KEYINPUT20), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  INV_X1    g094(.A(new_n282_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n266_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n278_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n243_), .B2(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n288_), .A2(new_n289_), .B1(new_n223_), .B2(new_n212_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n273_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n292_), .A2(new_n294_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n202_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT98), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n259_), .A2(new_n272_), .A3(KEYINPUT97), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT97), .B1(new_n259_), .B2(new_n272_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n243_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n300_), .B2(new_n283_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n294_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n295_), .B1(new_n300_), .B2(new_n283_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n294_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n274_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n308_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n310_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AOI211_X1 g120(.A(KEYINPUT98), .B(new_n308_), .C1(new_n315_), .C2(new_n318_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n309_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n316_), .B2(new_n274_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n317_), .B1(new_n243_), .B2(new_n273_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(new_n314_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n320_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n243_), .B2(new_n298_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n300_), .A2(new_n301_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n294_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n299_), .A2(new_n302_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n330_), .A2(KEYINPUT92), .A3(new_n308_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT92), .B1(new_n303_), .B2(new_n308_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n202_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n339_), .A2(new_n342_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(KEYINPUT1), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G155gat), .A3(G162gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n351_), .A3(new_n346_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G141gat), .B(G148gat), .Z(new_n353_));
  AOI22_X1  g152(.A1(new_n345_), .A2(new_n348_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT28), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n345_), .A2(new_n348_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n353_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n243_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n357_), .A2(new_n243_), .A3(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(G78gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G106gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n364_), .A2(new_n365_), .A3(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT93), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379_));
  INV_X1    g178(.A(G134gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G127gat), .ZN(new_n381_));
  INV_X1    g180(.A(G127gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G134gat), .ZN(new_n383_));
  INV_X1    g182(.A(G120gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G113gat), .ZN(new_n385_));
  INV_X1    g184(.A(G113gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G120gat), .ZN(new_n387_));
  AND4_X1   g186(.A1(new_n381_), .A2(new_n383_), .A3(new_n385_), .A4(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n381_), .A2(new_n383_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n379_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n379_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n361_), .A2(new_n390_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n391_), .B(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n354_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n396_), .B2(new_n379_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT4), .B1(new_n399_), .B2(new_n361_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n377_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n397_), .A3(new_n376_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n401_), .A2(new_n402_), .A3(new_n408_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n375_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n323_), .A2(new_n335_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n330_), .A2(new_n308_), .A3(new_n331_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(KEYINPUT33), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n401_), .A2(new_n420_), .A3(new_n402_), .A4(new_n408_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n395_), .A2(new_n397_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT95), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n395_), .A2(KEYINPUT95), .A3(new_n397_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n377_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n376_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n409_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT96), .B1(new_n418_), .B2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n327_), .A2(new_n332_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n429_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .A4(new_n417_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n319_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n303_), .A2(new_n437_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n439_), .A2(new_n412_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n431_), .A2(new_n436_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n414_), .B1(new_n443_), .B2(new_n375_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(KEYINPUT82), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G15gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT30), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n283_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n446_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n451_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT99), .B1(new_n444_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT99), .ZN(new_n457_));
  INV_X1    g256(.A(new_n375_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n432_), .A2(new_n434_), .A3(new_n417_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n441_), .B1(new_n459_), .B2(KEYINPUT96), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n460_), .B2(new_n436_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n457_), .B(new_n454_), .C1(new_n461_), .C2(new_n414_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n323_), .A2(new_n335_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n458_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n454_), .A2(new_n412_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT64), .B(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G85gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n474_), .B(KEYINPUT65), .Z(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT10), .B(G99gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n482_), .A2(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(KEYINPUT67), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n369_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n493_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G85gat), .B(G92gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n487_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AOI211_X1 g297(.A(new_n496_), .B(new_n486_), .C1(new_n490_), .C2(new_n494_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n484_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G57gat), .B(G64gat), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n503_));
  XOR2_X1   g302(.A(G71gat), .B(G78gat), .Z(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n503_), .A2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n500_), .A2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n484_), .B(new_n507_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(KEYINPUT12), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n500_), .A2(new_n512_), .A3(new_n508_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n469_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n468_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G120gat), .B(G148gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G176gat), .B(G204gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n514_), .A2(new_n515_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT13), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT13), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT75), .B(G1gat), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G8gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G29gat), .B(G36gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(KEYINPUT15), .A3(new_n542_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(new_n534_), .A3(new_n535_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT76), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n534_), .A2(new_n542_), .A3(new_n541_), .A4(new_n535_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n544_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n549_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n544_), .A2(new_n548_), .A3(new_n556_), .A4(new_n549_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT77), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT78), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n550_), .A2(KEYINPUT76), .B1(new_n553_), .B2(new_n554_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n565_), .A2(KEYINPUT78), .A3(new_n557_), .A4(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n557_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n561_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n507_), .B(new_n572_), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n536_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT17), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(KEYINPUT17), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n574_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n574_), .A2(new_n580_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n526_), .A2(new_n571_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT69), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n484_), .B(new_n543_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n495_), .A2(new_n497_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n486_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n495_), .A2(new_n497_), .A3(new_n487_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n483_), .A2(new_n481_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n597_), .A2(new_n598_), .B1(new_n476_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n546_), .A2(new_n547_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n590_), .B(new_n595_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT72), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n589_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n500_), .A2(new_n547_), .A3(new_n546_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(KEYINPUT69), .A3(new_n590_), .A4(new_n595_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n593_), .A2(new_n594_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  OAI221_X1 g407(.A(new_n589_), .B1(new_n594_), .B2(new_n593_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(KEYINPUT73), .A3(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n609_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n616_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n610_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n610_), .B1(new_n619_), .B2(new_n618_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n587_), .B(new_n588_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n608_), .A2(new_n609_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n619_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n623_), .B(KEYINPUT73), .C1(new_n624_), .C2(new_n617_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n610_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(KEYINPUT74), .A3(new_n586_), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n585_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n467_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT100), .Z(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n412_), .A3(new_n527_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n625_), .A2(new_n626_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n467_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n585_), .B(KEYINPUT101), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n412_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n633_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  NAND3_X1  g442(.A1(new_n631_), .A2(new_n528_), .A3(new_n463_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n637_), .A2(new_n463_), .A3(new_n638_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n528_), .B1(new_n645_), .B2(KEYINPUT102), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n637_), .A2(new_n638_), .A3(new_n648_), .A4(new_n463_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n644_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT40), .B(new_n644_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n639_), .B2(new_n454_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n658_), .ZN(new_n660_));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n631_), .A2(new_n661_), .A3(new_n455_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n639_), .B2(new_n375_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n631_), .A2(new_n667_), .A3(new_n458_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n584_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n526_), .A2(new_n571_), .A3(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n636_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n467_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n467_), .A2(new_n672_), .A3(KEYINPUT106), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n412_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n467_), .A2(new_n628_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n467_), .A2(new_n681_), .A3(new_n628_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n671_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT105), .B1(new_n683_), .B2(KEYINPUT44), .ZN(new_n684_));
  INV_X1    g483(.A(new_n671_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n467_), .A2(new_n681_), .A3(new_n628_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n681_), .B1(new_n467_), .B2(new_n628_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n685_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(G29gat), .A3(new_n412_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n678_), .B1(new_n692_), .B2(new_n694_), .ZN(G1328gat));
  XOR2_X1   g494(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n696_));
  INV_X1    g495(.A(new_n463_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n677_), .B2(new_n698_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n675_), .A2(new_n676_), .A3(new_n696_), .A4(new_n698_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n693_), .A2(new_n463_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n684_), .B2(new_n691_), .ZN(new_n703_));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  OAI221_X1 g507(.A(new_n701_), .B1(new_n706_), .B2(KEYINPUT46), .C1(new_n703_), .C2(new_n704_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n693_), .A2(G43gat), .A3(new_n455_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n684_), .B2(new_n691_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G43gat), .B1(new_n677_), .B2(new_n455_), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n712_), .A2(new_n713_), .A3(KEYINPUT47), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT47), .B1(new_n712_), .B2(new_n713_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n677_), .B2(new_n458_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n693_), .A2(G50gat), .A3(new_n458_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n692_), .B2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(new_n571_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n526_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n720_), .A2(new_n637_), .A3(new_n721_), .A4(new_n584_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n412_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G57gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n467_), .A2(new_n720_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n526_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n628_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n467_), .A2(KEYINPUT109), .A3(new_n720_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n727_), .A2(new_n584_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n640_), .A2(G57gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n724_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g532(.A(G64gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n722_), .B2(new_n463_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT48), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n463_), .A2(new_n734_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n730_), .B2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n722_), .B2(new_n455_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT49), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n455_), .A2(new_n739_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n730_), .B2(new_n742_), .ZN(G1334gat));
  AOI21_X1  g542(.A(new_n367_), .B1(new_n722_), .B2(new_n458_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT50), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n458_), .A2(new_n367_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n730_), .B2(new_n746_), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n636_), .A2(new_n584_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n727_), .A2(new_n729_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT111), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n727_), .A2(new_n751_), .A3(new_n729_), .A4(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(G85gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n412_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n680_), .A2(new_n682_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n526_), .A2(new_n571_), .A3(new_n584_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n412_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n754_), .B2(new_n760_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n463_), .A3(new_n470_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n697_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G92gat), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n762_), .B(KEYINPUT112), .C1(new_n763_), .C2(G92gat), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1337gat));
  OAI211_X1 g567(.A(new_n455_), .B(new_n757_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G99gat), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT113), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n454_), .B(new_n482_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n770_), .B(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n454_), .A2(new_n482_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n753_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(new_n779_), .ZN(G1338gat));
  OAI211_X1 g579(.A(new_n458_), .B(new_n757_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G106gat), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n782_), .B(new_n784_), .ZN(new_n785_));
  AOI211_X1 g584(.A(G106gat), .B(new_n375_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT53), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n782_), .B(new_n783_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n753_), .A2(new_n369_), .A3(new_n458_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(G1339gat));
  NAND3_X1  g591(.A1(new_n464_), .A2(new_n455_), .A3(new_n412_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n511_), .A2(new_n513_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n468_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n514_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n514_), .A2(new_n797_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n520_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n794_), .B(KEYINPUT56), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n553_), .A2(new_n549_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n544_), .A2(new_n548_), .A3(new_n554_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n569_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n567_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT116), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n567_), .A2(new_n808_), .A3(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n514_), .A2(new_n797_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT55), .B(new_n469_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n812_));
  OAI22_X1  g611(.A1(new_n811_), .A2(new_n812_), .B1(new_n468_), .B2(new_n795_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT119), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n794_), .A2(KEYINPUT56), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n813_), .A2(new_n520_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n802_), .A2(new_n810_), .A3(new_n521_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n514_), .A2(new_n515_), .A3(new_n520_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n822_), .A2(new_n802_), .A3(KEYINPUT58), .A4(new_n817_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n628_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n820_), .A2(new_n628_), .A3(KEYINPUT120), .A4(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n800_), .A2(new_n801_), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n813_), .A2(new_n830_), .A3(new_n814_), .A4(new_n520_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n821_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n521_), .A2(new_n522_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n809_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n808_), .B1(new_n567_), .B2(new_n805_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n635_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n839_), .B2(KEYINPUT57), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n831_), .A2(new_n832_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n813_), .A2(new_n520_), .B1(new_n830_), .B2(new_n814_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n636_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n839_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n841_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n670_), .B1(new_n828_), .B2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n728_), .A2(new_n720_), .A3(new_n526_), .A4(new_n584_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT54), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n793_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853_), .B2(new_n571_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n793_), .A2(KEYINPUT59), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT118), .B1(new_n838_), .B2(new_n845_), .ZN(new_n858_));
  OAI22_X1  g657(.A1(new_n858_), .A2(KEYINPUT57), .B1(new_n838_), .B2(new_n840_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n584_), .B1(new_n859_), .B2(new_n824_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n851_), .B(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n857_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n386_), .B1(new_n571_), .B2(KEYINPUT121), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(KEYINPUT121), .B2(new_n386_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n854_), .B1(new_n865_), .B2(new_n867_), .ZN(G1340gat));
  OAI211_X1 g667(.A(new_n863_), .B(new_n721_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n384_), .B1(new_n526_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n853_), .B(new_n871_), .C1(KEYINPUT60), .C2(new_n384_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(KEYINPUT122), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n864_), .B2(new_n670_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n853_), .A2(new_n382_), .A3(new_n584_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n853_), .B2(new_n635_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT123), .B(G134gat), .Z(new_n882_));
  NOR2_X1   g681(.A1(new_n728_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n865_), .B2(new_n883_), .ZN(G1343gat));
  AOI21_X1  g683(.A(new_n455_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n463_), .A2(new_n640_), .A3(new_n375_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n720_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n337_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n526_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n338_), .ZN(G1345gat));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n670_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n892_), .B(new_n893_), .Z(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n887_), .B2(new_n728_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n636_), .A2(G162gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n887_), .B2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n860_), .A2(new_n862_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n465_), .A2(new_n463_), .A3(new_n375_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n720_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n898_), .B(new_n899_), .C1(new_n903_), .C2(new_n261_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n261_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n905_));
  OAI221_X1 g704(.A(new_n905_), .B1(KEYINPUT124), .B2(KEYINPUT62), .C1(new_n902_), .C2(new_n720_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n256_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  INV_X1    g707(.A(new_n902_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G176gat), .B1(new_n909_), .B2(new_n721_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n901_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(G176gat), .A3(new_n721_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n910_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n670_), .A2(new_n267_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n909_), .B2(new_n917_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n902_), .A2(KEYINPUT126), .A3(new_n267_), .A4(new_n670_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n911_), .B2(new_n584_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n902_), .B2(new_n728_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n635_), .A2(new_n268_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n902_), .B2(new_n923_), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n463_), .A2(new_n413_), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n455_), .B(new_n925_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(G197gat), .A3(new_n571_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G197gat), .B1(new_n926_), .B2(new_n571_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n926_), .A2(new_n721_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g733(.A(KEYINPUT63), .B(G211gat), .C1(new_n926_), .C2(new_n584_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n926_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n670_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AOI21_X1  g737(.A(new_n935_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n936_), .B2(new_n728_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n926_), .A2(new_n203_), .A3(new_n635_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1355gat));
endmodule


