//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT34), .Z(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G85gat), .B(G92gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT8), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT65), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT7), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n208_), .B1(KEYINPUT65), .B2(new_n210_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n207_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n218_), .B2(new_n220_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n227_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n206_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT67), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT67), .B1(new_n228_), .B2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n222_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234_));
  INV_X1    g033(.A(G92gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n206_), .B1(KEYINPUT9), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(KEYINPUT9), .B2(new_n206_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(KEYINPUT64), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(KEYINPUT64), .ZN(new_n239_));
  INV_X1    g038(.A(G106gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT10), .B(G99gat), .Z(new_n241_));
  AOI21_X1  g040(.A(new_n221_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n233_), .A2(new_n234_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n234_), .B1(new_n233_), .B2(new_n243_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G29gat), .B(G36gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT73), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n244_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n203_), .A2(new_n204_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT74), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(KEYINPUT75), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n233_), .A2(new_n243_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n251_), .B(KEYINPUT15), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n255_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n205_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G190gat), .B(G218gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G134gat), .B(G162gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT36), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n256_), .A2(KEYINPUT68), .ZN(new_n265_));
  INV_X1    g064(.A(new_n251_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n233_), .A2(new_n234_), .A3(new_n243_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n205_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT15), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n251_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n256_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n268_), .A2(new_n269_), .A3(new_n272_), .A4(new_n255_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n260_), .A2(new_n264_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n260_), .A2(new_n273_), .A3(KEYINPUT76), .A4(new_n264_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n260_), .A2(new_n273_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n263_), .B(KEYINPUT36), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT77), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT37), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT37), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n284_), .A3(new_n274_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n281_), .B2(KEYINPUT37), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT78), .B(G15gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G22gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G71gat), .B(G78gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n300_), .B(new_n308_), .Z(new_n309_));
  XOR2_X1   g108(.A(G127gat), .B(G155gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT16), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G183gat), .B(G211gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT17), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT79), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n313_), .A2(new_n314_), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n309_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n288_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G229gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n271_), .A2(new_n298_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT80), .B1(new_n298_), .B2(new_n251_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n266_), .A2(new_n326_), .A3(new_n297_), .A4(new_n296_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n323_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G169gat), .B(G197gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(KEYINPUT81), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n298_), .A2(new_n251_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n334_), .C1(new_n322_), .C2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n322_), .ZN(new_n338_));
  OAI22_X1  g137(.A1(new_n338_), .A2(new_n329_), .B1(KEYINPUT81), .B2(new_n333_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT82), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(G183gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G183gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(KEYINPUT25), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT84), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n347_), .B2(KEYINPUT25), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n346_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT23), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(G183gat), .A3(G190gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n356_), .A2(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT85), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n361_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G169gat), .ZN(new_n366_));
  INV_X1    g165(.A(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n362_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n355_), .A2(new_n357_), .ZN(new_n371_));
  INV_X1    g170(.A(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n347_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n368_), .B(new_n370_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n358_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT86), .B1(new_n378_), .B2(new_n373_), .ZN(new_n379_));
  OAI22_X1  g178(.A1(new_n354_), .A2(new_n365_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT87), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n384_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(G15gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n387_), .A2(new_n391_), .ZN(new_n394_));
  OR3_X1    g193(.A1(new_n393_), .A2(KEYINPUT88), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT88), .B1(new_n393_), .B2(new_n394_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  OAI211_X1 g201(.A(KEYINPUT88), .B(new_n402_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(KEYINPUT97), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n411_));
  AND2_X1   g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT95), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n344_), .A2(new_n348_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n364_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n417_), .A2(new_n350_), .B1(new_n362_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n361_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n360_), .A2(new_n359_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n378_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n368_), .A2(new_n370_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n375_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G197gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G204gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT21), .ZN(new_n433_));
  INV_X1    g232(.A(G204gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G197gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .A4(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G211gat), .B(G218gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n433_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT91), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n440_));
  AOI211_X1 g239(.A(new_n440_), .B(new_n433_), .C1(new_n429_), .C2(new_n435_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n436_), .B(new_n437_), .C1(new_n439_), .C2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n437_), .A2(new_n433_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n431_), .A2(new_n435_), .A3(new_n432_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n416_), .B1(new_n427_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n438_), .B(KEYINPUT91), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n436_), .A2(new_n437_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n448_), .A2(new_n449_), .B1(new_n444_), .B2(new_n443_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n377_), .A2(new_n379_), .ZN(new_n451_));
  OAI221_X1 g250(.A(new_n361_), .B1(new_n363_), .B2(new_n364_), .C1(new_n346_), .C2(new_n353_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n415_), .B1(new_n447_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n427_), .B2(new_n446_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n380_), .A2(new_n446_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n410_), .A2(new_n454_), .B1(new_n457_), .B2(new_n413_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n447_), .A2(new_n453_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n414_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT97), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n409_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n361_), .B(new_n420_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n463_), .A2(new_n419_), .B1(new_n425_), .B2(new_n375_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n464_), .B2(new_n450_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n380_), .A2(new_n446_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n410_), .B(new_n414_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n416_), .B1(new_n464_), .B2(new_n450_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n468_), .B(new_n413_), .C1(new_n450_), .C2(new_n381_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n409_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n410_), .B1(new_n459_), .B2(new_n414_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n405_), .B1(new_n462_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n458_), .A2(new_n409_), .A3(new_n461_), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n457_), .A2(new_n413_), .B1(new_n459_), .B2(new_n414_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n405_), .B1(new_n476_), .B2(new_n471_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n477_), .A3(KEYINPUT101), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT101), .B1(new_n475_), .B2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n474_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G141gat), .A2(G148gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT89), .ZN(new_n483_));
  AND2_X1   g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n484_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n483_), .B(new_n485_), .C1(KEYINPUT1), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G141gat), .A2(G148gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT2), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n491_), .A2(new_n494_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n487_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n489_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT29), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n446_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G228gat), .A2(G233gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT90), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n502_), .B(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT28), .B1(new_n499_), .B2(KEYINPUT29), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n489_), .A2(new_n508_), .A3(new_n501_), .A4(new_n498_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G22gat), .B(G50gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n506_), .B(KEYINPUT93), .C1(new_n512_), .C2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT93), .B1(new_n512_), .B2(new_n513_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n513_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n511_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n502_), .B(new_n504_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G78gat), .B(G106gat), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n514_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G29gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G85gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT4), .ZN(new_n534_));
  INV_X1    g333(.A(new_n399_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n500_), .A2(KEYINPUT98), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n499_), .A2(new_n399_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(KEYINPUT98), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n534_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(KEYINPUT4), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n533_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(new_n540_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(new_n533_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n531_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n531_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n481_), .A2(new_n526_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n524_), .A2(new_n525_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n458_), .A2(new_n461_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(KEYINPUT100), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n476_), .A2(new_n554_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT100), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n551_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n462_), .A2(new_n473_), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT33), .B(new_n531_), .C1(new_n544_), .C2(new_n546_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n549_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n541_), .A2(new_n533_), .A3(new_n542_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n531_), .B1(new_n545_), .B2(new_n533_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n562_), .B(new_n563_), .C1(new_n564_), .C2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n553_), .B1(new_n561_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n404_), .B1(new_n552_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n404_), .A2(new_n551_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT102), .ZN(new_n573_));
  INV_X1    g372(.A(new_n480_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n478_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n573_), .B1(new_n575_), .B2(new_n474_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n474_), .B(new_n573_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n526_), .B(new_n572_), .C1(new_n576_), .C2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n342_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n244_), .A2(new_n245_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n308_), .ZN(new_n584_));
  INV_X1    g383(.A(G230gat), .ZN(new_n585_));
  INV_X1    g384(.A(G233gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n583_), .B2(new_n308_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n256_), .A2(KEYINPUT12), .A3(new_n307_), .A4(new_n306_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n265_), .A2(new_n308_), .A3(new_n267_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n308_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n587_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G120gat), .B(G148gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n590_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n603_));
  AND2_X1   g402(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n604_));
  NOR2_X1   g403(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n602_), .B(new_n603_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n602_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n603_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n609_), .B2(new_n605_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n321_), .A2(new_n580_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n551_), .B(KEYINPUT103), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n612_), .A2(new_n291_), .A3(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n340_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n320_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n280_), .A2(new_n620_), .A3(new_n274_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n280_), .B2(new_n274_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n551_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n615_), .A2(new_n616_), .A3(new_n627_), .ZN(G1324gat));
  NOR2_X1   g427(.A1(new_n576_), .A2(new_n578_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n612_), .A2(new_n292_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G8gat), .B1(new_n625_), .B2(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT105), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(KEYINPUT105), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n630_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT40), .B(new_n630_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1325gat));
  OAI21_X1  g441(.A(G15gat), .B1(new_n625_), .B2(new_n404_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n611_), .A2(G15gat), .A3(new_n404_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(G1326gat));
  OAI21_X1  g447(.A(G22gat), .B1(new_n625_), .B2(new_n526_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n526_), .A2(G22gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n611_), .B2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(G29gat), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n571_), .A2(new_n579_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n281_), .A2(KEYINPUT37), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT77), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n658_), .A2(KEYINPUT107), .A3(new_n285_), .A4(new_n283_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT43), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT43), .B1(new_n571_), .B2(new_n579_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n288_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(KEYINPUT44), .A3(new_n320_), .A4(new_n618_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n660_), .A2(KEYINPUT43), .B1(new_n288_), .B2(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n618_), .A2(new_n320_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n653_), .B1(new_n670_), .B2(new_n613_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n623_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n619_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n580_), .A2(new_n610_), .A3(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(G29gat), .A3(new_n626_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n671_), .A2(new_n675_), .ZN(G1328gat));
  OR2_X1    g475(.A1(new_n629_), .A2(KEYINPUT109), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n629_), .A2(KEYINPUT109), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n674_), .A2(G36gat), .A3(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT45), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n665_), .A2(new_n669_), .A3(new_n629_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G36gat), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT46), .B(new_n681_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  NOR3_X1   g489(.A1(new_n674_), .A2(G43gat), .A3(new_n404_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n404_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n665_), .A2(new_n669_), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n693_), .B2(G43gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n670_), .A2(new_n553_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(G50gat), .ZN(new_n698_));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT110), .B(new_n699_), .C1(new_n670_), .C2(new_n553_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n553_), .A2(new_n699_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n698_), .A2(new_n700_), .B1(new_n674_), .B2(new_n701_), .ZN(G1331gat));
  AOI211_X1 g501(.A(new_n340_), .B(new_n610_), .C1(new_n571_), .C2(new_n579_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n321_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT111), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT111), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n613_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G57gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n610_), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n342_), .A2(new_n624_), .A3(new_n710_), .A4(new_n619_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n626_), .A2(new_n709_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n708_), .A2(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n679_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n705_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n711_), .B2(new_n692_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT49), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n705_), .A2(new_n720_), .A3(new_n692_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n711_), .B2(new_n553_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT50), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n705_), .A2(new_n725_), .A3(new_n553_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1335gat));
  AND2_X1   g528(.A1(new_n703_), .A2(new_n673_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n613_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(G85gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT112), .Z(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n661_), .A2(new_n735_), .A3(new_n663_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n610_), .A2(new_n340_), .A3(new_n619_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n667_), .A2(new_n735_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n664_), .A2(KEYINPUT113), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT114), .A3(new_n737_), .A4(new_n736_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n740_), .A2(new_n742_), .A3(G85gat), .A4(new_n551_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n733_), .A2(new_n743_), .ZN(G1336gat));
  NAND3_X1  g543(.A1(new_n730_), .A2(new_n235_), .A3(new_n629_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n740_), .A2(new_n715_), .A3(new_n742_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n235_), .ZN(G1337gat));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n692_), .A3(new_n742_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(G99gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n730_), .A2(new_n692_), .A3(new_n241_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT51), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n753_), .A3(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1338gat));
  AND2_X1   g554(.A1(new_n737_), .A2(new_n553_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n240_), .B1(new_n664_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n730_), .A2(new_n240_), .A3(new_n553_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n589_), .B1(new_n593_), .B2(new_n581_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n591_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n584_), .A2(new_n588_), .A3(KEYINPUT55), .A4(new_n589_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n591_), .B(new_n589_), .C1(new_n593_), .C2(new_n581_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n587_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n601_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT115), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n771_), .A2(KEYINPUT115), .A3(new_n773_), .A4(new_n601_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n340_), .A2(new_n603_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n333_), .B1(new_n338_), .B2(new_n329_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n336_), .A2(new_n323_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n324_), .A2(new_n328_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n323_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n783_), .B2(new_n333_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n623_), .B1(new_n779_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n763_), .B1(new_n787_), .B2(KEYINPUT57), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n777_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n790_), .B2(new_n776_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT116), .B(new_n789_), .C1(new_n791_), .C2(new_n623_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n787_), .A2(KEYINPUT57), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n608_), .A2(new_n784_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n771_), .A2(new_n773_), .A3(new_n601_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n773_), .B1(new_n771_), .B2(new_n601_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n798_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n800_), .A2(KEYINPUT58), .A3(new_n796_), .A4(new_n795_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n288_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n788_), .A2(new_n792_), .A3(new_n793_), .A4(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n658_), .A2(new_n285_), .A3(new_n283_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n610_), .A3(new_n619_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT54), .B1(new_n805_), .B2(new_n341_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n321_), .A2(new_n807_), .A3(new_n342_), .A4(new_n610_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n803_), .A2(new_n320_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n629_), .A2(new_n553_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n692_), .A3(new_n613_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n340_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n803_), .A2(new_n320_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n808_), .A2(new_n806_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n811_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n793_), .A2(new_n802_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n787_), .A2(KEYINPUT57), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n320_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n815_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n817_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n819_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT117), .B(G113gat), .Z(new_n828_));
  NAND2_X1  g627(.A1(new_n341_), .A2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT118), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n813_), .B1(new_n827_), .B2(new_n830_), .ZN(G1340gat));
  OAI211_X1 g630(.A(new_n710_), .B(new_n825_), .C1(new_n812_), .C2(new_n824_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT119), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n819_), .A2(new_n834_), .A3(new_n710_), .A4(new_n825_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n835_), .A3(G120gat), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n812_), .B(new_n838_), .C1(KEYINPUT60), .C2(new_n837_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1341gat));
  NAND2_X1  g639(.A1(new_n619_), .A2(G127gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT120), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n825_), .B(new_n842_), .C1(new_n812_), .C2(new_n824_), .ZN(new_n843_));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n818_), .B2(new_n320_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT121), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n845_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1342gat));
  OAI21_X1  g649(.A(G134gat), .B1(new_n826_), .B2(new_n804_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n672_), .A2(G134gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n818_), .B2(new_n852_), .ZN(G1343gat));
  NAND3_X1  g652(.A1(new_n679_), .A2(new_n553_), .A3(new_n613_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n809_), .A2(new_n692_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n340_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n710_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n619_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  AOI21_X1  g661(.A(G162gat), .B1(new_n855_), .B2(new_n623_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n655_), .A2(G162gat), .A3(new_n659_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n855_), .B2(new_n864_), .ZN(G1347gat));
  INV_X1    g664(.A(G169gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n613_), .A2(new_n404_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n715_), .A2(new_n526_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n822_), .B2(new_n815_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n340_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT123), .ZN(new_n873_));
  INV_X1    g672(.A(new_n871_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n869_), .A2(new_n340_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT124), .B(new_n874_), .C1(new_n875_), .C2(new_n866_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n870_), .A2(new_n879_), .A3(new_n871_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n873_), .A2(new_n876_), .A3(new_n878_), .A4(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n875_), .A2(new_n366_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(G176gat), .B1(new_n869_), .B2(new_n710_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n809_), .A2(new_n553_), .ZN(new_n885_));
  AND4_X1   g684(.A1(G176gat), .A2(new_n710_), .A3(new_n715_), .A4(new_n867_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  INV_X1    g686(.A(new_n868_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n823_), .A2(new_n888_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n889_), .A2(new_n417_), .A3(new_n320_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n885_), .A2(new_n619_), .A3(new_n715_), .A4(new_n867_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n347_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n889_), .B2(new_n804_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n869_), .A2(new_n350_), .A3(new_n623_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1351gat));
  XNOR2_X1  g696(.A(KEYINPUT127), .B(G197gat), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n679_), .A2(new_n551_), .A3(new_n526_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n816_), .A2(new_n404_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT126), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n692_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n899_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n898_), .B1(new_n905_), .B2(new_n340_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n428_), .A2(KEYINPUT127), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n903_), .B1(new_n902_), .B2(new_n899_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n899_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n809_), .A2(KEYINPUT126), .A3(new_n692_), .A4(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n340_), .B(new_n907_), .C1(new_n908_), .C2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n906_), .A2(new_n912_), .ZN(G1352gat));
  OAI21_X1  g712(.A(new_n710_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n905_), .B2(new_n619_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT63), .B(G211gat), .Z(new_n918_));
  OAI211_X1 g717(.A(new_n619_), .B(new_n918_), .C1(new_n908_), .C2(new_n910_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n920_), .ZN(G1354gat));
  INV_X1    g720(.A(G218gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n905_), .A2(new_n922_), .A3(new_n623_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n804_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1355gat));
endmodule


