//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n972_, new_n973_, new_n974_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  AND3_X1   g003(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT1), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT84), .ZN(new_n214_));
  INV_X1    g013(.A(G155gat), .ZN(new_n215_));
  INV_X1    g014(.A(G162gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n207_), .A2(new_n213_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n218_), .A2(new_n217_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n204_), .B1(new_n225_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n220_), .A2(new_n224_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n204_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G225gat), .A2(G233gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT92), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n225_), .A2(new_n234_), .A3(new_n204_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n243_), .A2(new_n235_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n225_), .A2(new_n234_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n204_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n240_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n242_), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G1gat), .B(G29gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G85gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n242_), .B(new_n255_), .C1(new_n245_), .C2(new_n250_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(G15gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT30), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT23), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT77), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G190gat), .ZN(new_n274_));
  INV_X1    g073(.A(G183gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n272_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n270_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT81), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n280_));
  NOR2_X1   g079(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n281_));
  OAI21_X1  g080(.A(G169gat), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT80), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(G169gat), .C1(new_n280_), .C2(new_n281_), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  AOI21_X1  g085(.A(G176gat), .B1(new_n286_), .B2(KEYINPUT22), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n267_), .A2(new_n289_), .A3(new_n276_), .A4(new_n270_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n278_), .A2(new_n279_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT78), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n268_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT23), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n269_), .B1(G183gat), .B2(G190gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n286_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n279_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(KEYINPUT24), .ZN(new_n302_));
  NOR2_X1   g101(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n272_), .A2(new_n274_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(KEYINPUT26), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n306_), .A2(new_n275_), .A3(KEYINPUT25), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(KEYINPUT25), .B2(new_n275_), .ZN(new_n308_));
  OAI22_X1  g107(.A1(new_n307_), .A2(new_n308_), .B1(KEYINPUT25), .B2(new_n275_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n297_), .B(new_n302_), .C1(new_n305_), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n291_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G71gat), .B(G99gat), .ZN(new_n312_));
  INV_X1    g111(.A(G43gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n311_), .A2(new_n314_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n264_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n311_), .A2(new_n314_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n263_), .A3(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT82), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  AOI211_X1 g124(.A(new_n324_), .B(new_n325_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n318_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT83), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n259_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n267_), .A2(new_n270_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT25), .B(G183gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n301_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(new_n299_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n286_), .A2(KEYINPUT22), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT22), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G169gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n348_), .A3(new_n298_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n279_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(KEYINPUT90), .A3(new_n279_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n275_), .A2(new_n271_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT91), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n349_), .A2(KEYINPUT90), .A3(new_n279_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT90), .B1(new_n349_), .B2(new_n279_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n356_), .B(KEYINPUT91), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n345_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G211gat), .B(G218gat), .Z(new_n363_));
  INV_X1    g162(.A(G197gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G204gat), .ZN(new_n365_));
  INV_X1    g164(.A(G204gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G197gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n363_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT87), .B1(new_n368_), .B2(KEYINPUT21), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT21), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n365_), .A2(new_n367_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT86), .B1(new_n366_), .B2(G197gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n364_), .A3(G204gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n377_), .A3(new_n367_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n363_), .B1(new_n378_), .B2(KEYINPUT21), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n369_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n362_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n291_), .A2(new_n310_), .A3(new_n380_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n337_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n360_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n380_), .A3(new_n345_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n337_), .A2(KEYINPUT20), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n311_), .B2(new_n381_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n334_), .B1(new_n385_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n380_), .B1(new_n389_), .B2(new_n345_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n383_), .A2(KEYINPUT20), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n336_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n334_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(new_n392_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  AND4_X1   g201(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n388_), .B2(new_n360_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT20), .B(new_n383_), .C1(new_n404_), .C2(new_n380_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n405_), .A2(new_n336_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n402_), .B1(new_n406_), .B2(new_n398_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n336_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n380_), .A2(new_n345_), .A3(new_n386_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n409_), .A2(KEYINPUT20), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n311_), .A2(new_n381_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n337_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n334_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n401_), .A2(new_n402_), .B1(new_n407_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n246_), .A2(KEYINPUT29), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n381_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n225_), .B2(new_n234_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n420_), .B2(new_n380_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n237_), .A2(new_n419_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT28), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n428_), .B(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n424_), .A2(new_n431_), .A3(new_n433_), .A4(new_n426_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT95), .B1(new_n414_), .B2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n398_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n402_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n413_), .A2(KEYINPUT27), .A3(new_n400_), .ZN(new_n442_));
  AND4_X1   g241(.A1(KEYINPUT95), .A2(new_n441_), .A3(new_n437_), .A4(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n330_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n328_), .B(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n323_), .A2(new_n326_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n435_), .A2(new_n436_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n259_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n441_), .A2(new_n442_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n258_), .B2(KEYINPUT94), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n249_), .A2(new_n241_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n245_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n236_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n256_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n258_), .A2(KEYINPUT94), .A3(new_n453_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n400_), .A3(new_n394_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n398_), .A2(KEYINPUT32), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n406_), .A2(new_n463_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n259_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n449_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n448_), .B1(new_n452_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n444_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT15), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT73), .B(G1gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n482_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n476_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n478_), .A2(new_n484_), .A3(new_n487_), .A4(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n484_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n476_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n477_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n471_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G141gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n470_), .A2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n502_), .A2(KEYINPUT96), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(KEYINPUT96), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G120gat), .B(G148gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT65), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(G85gat), .A3(G92gat), .A4(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n515_), .A2(new_n511_), .A3(KEYINPUT9), .A4(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT6), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n527_), .A3(KEYINPUT66), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n535_));
  INV_X1    g334(.A(G99gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n519_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n530_), .A2(new_n531_), .A3(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n515_), .A2(new_n516_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n525_), .A2(new_n527_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n537_), .A2(new_n538_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n541_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT8), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n544_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n534_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(KEYINPUT11), .B2(new_n553_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT12), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n552_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT64), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n540_), .A2(new_n543_), .B1(new_n548_), .B2(KEYINPUT8), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n522_), .A2(new_n532_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n560_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n566_), .A2(new_n560_), .A3(new_n567_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n565_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n544_), .A2(new_n549_), .B1(new_n523_), .B2(new_n533_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n559_), .A2(new_n558_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n573_), .B1(new_n577_), .B2(new_n569_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n510_), .B1(new_n572_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n578_), .A3(new_n510_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n572_), .A2(new_n578_), .A3(new_n510_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n584_), .A2(new_n579_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT69), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n544_), .A2(new_n549_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n476_), .A3(new_n534_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n478_), .A2(new_n489_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n599_), .B2(new_n552_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n594_), .A2(new_n595_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n589_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n574_), .A2(new_n476_), .B1(new_n595_), .B2(new_n594_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n590_), .A2(KEYINPUT67), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n566_), .A2(new_n545_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n567_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n607_), .B2(new_n598_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(KEYINPUT69), .A3(new_n601_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n603_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n600_), .A2(KEYINPUT71), .A3(new_n602_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n602_), .B(new_n604_), .C1(new_n607_), .C2(new_n598_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT71), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT70), .ZN(new_n617_));
  XOR2_X1   g416(.A(G134gat), .B(G162gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n610_), .A2(new_n615_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT72), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n588_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n603_), .A2(new_n609_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n619_), .B(KEYINPUT36), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  OAI221_X1 g429(.A(new_n623_), .B1(new_n624_), .B2(new_n588_), .C1(new_n626_), .C2(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n576_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(new_n491_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT74), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT16), .ZN(new_n639_));
  XOR2_X1   g438(.A(G183gat), .B(G211gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT17), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n637_), .B(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n635_), .A2(KEYINPUT17), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n632_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n505_), .A2(new_n587_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n259_), .A3(new_n479_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n450_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n441_), .A2(new_n442_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n449_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n414_), .A2(KEYINPUT95), .A3(new_n437_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n327_), .A2(new_n329_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n454_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n459_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n461_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n467_), .B1(new_n661_), .B2(new_n401_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n437_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n663_), .B2(new_n451_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n657_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n629_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n586_), .A2(new_n501_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT97), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(new_n646_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G1gat), .B1(new_n671_), .B2(new_n450_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n649_), .A2(new_n650_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n651_), .A2(new_n672_), .A3(new_n673_), .ZN(G1324gat));
  NAND3_X1  g473(.A1(new_n648_), .A2(new_n480_), .A3(new_n654_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n670_), .A2(new_n654_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G8gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT39), .B(new_n480_), .C1(new_n670_), .C2(new_n654_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1325gat));
  AND3_X1   g481(.A1(new_n648_), .A2(new_n261_), .A3(new_n658_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT100), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n670_), .A2(new_n658_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G15gat), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT99), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT41), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(KEYINPUT41), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n684_), .A2(new_n688_), .A3(new_n689_), .ZN(G1326gat));
  INV_X1    g489(.A(G22gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n670_), .B2(new_n449_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT42), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n648_), .A2(new_n691_), .A3(new_n449_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1327gat));
  INV_X1    g494(.A(new_n646_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n666_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n505_), .A2(new_n587_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n259_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n630_), .A2(new_n631_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n470_), .A2(KEYINPUT102), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT102), .B1(new_n470_), .B2(new_n704_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(new_n657_), .B2(new_n664_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n444_), .A2(new_n469_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n632_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT43), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n707_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n669_), .A2(new_n696_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n701_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT103), .B(new_n715_), .C1(new_n707_), .C2(new_n713_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n700_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n259_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n699_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n632_), .B1(new_n470_), .B2(KEYINPUT101), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n702_), .B1(new_n728_), .B2(new_n710_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n665_), .B2(new_n703_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n470_), .A2(new_n704_), .A3(KEYINPUT102), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n716_), .B1(new_n729_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n414_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n727_), .B1(new_n719_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n697_), .A2(new_n587_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n414_), .A2(G36gat), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n739_), .B(new_n740_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT45), .Z(new_n742_));
  OAI21_X1  g541(.A(new_n726_), .B1(new_n738_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n700_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n734_), .A2(KEYINPUT103), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n714_), .A2(new_n701_), .A3(new_n716_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n720_), .A2(new_n654_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G36gat), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n726_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n742_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n743_), .A2(new_n752_), .ZN(G1329gat));
  NAND2_X1  g552(.A1(new_n658_), .A2(G43gat), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n747_), .A2(new_n736_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G43gat), .B1(new_n698_), .B2(new_n658_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT47), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n758_));
  INV_X1    g557(.A(new_n756_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n758_), .B(new_n759_), .C1(new_n721_), .C2(new_n754_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1330gat));
  AOI21_X1  g560(.A(G50gat), .B1(new_n698_), .B2(new_n449_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n449_), .A2(G50gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n722_), .B2(new_n763_), .ZN(G1331gat));
  INV_X1    g563(.A(new_n500_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n497_), .B(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n470_), .A2(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(new_n586_), .A3(new_n647_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT106), .Z(new_n769_));
  INV_X1    g568(.A(G57gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n259_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n667_), .A2(new_n766_), .A3(new_n587_), .A4(new_n646_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G57gat), .B1(new_n772_), .B2(new_n450_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1332gat));
  INV_X1    g573(.A(G64gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n769_), .A2(new_n775_), .A3(new_n654_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G64gat), .B1(new_n772_), .B2(new_n414_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT48), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n772_), .B2(new_n448_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT107), .Z(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT49), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT49), .ZN(new_n783_));
  INV_X1    g582(.A(G71gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n769_), .A2(new_n784_), .A3(new_n658_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n769_), .A2(new_n787_), .A3(new_n449_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G78gat), .B1(new_n772_), .B2(new_n437_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT50), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1335gat));
  OR3_X1    g590(.A1(new_n767_), .A2(new_n586_), .A3(new_n697_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n792_), .A2(G85gat), .A3(new_n450_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n646_), .A2(new_n586_), .A3(new_n501_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n714_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n259_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n796_), .B2(G85gat), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(G1336gat));
  INV_X1    g598(.A(new_n792_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G92gat), .B1(new_n800_), .B2(new_n654_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n654_), .A2(G92gat), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT109), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n795_), .B2(new_n803_), .ZN(G1337gat));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n658_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n792_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n795_), .A2(new_n658_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(G99gat), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1338gat));
  NAND3_X1  g610(.A1(new_n800_), .A2(new_n519_), .A3(new_n449_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n714_), .A2(new_n449_), .A3(new_n794_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815_));
  AND4_X1   g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .A4(G106gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n519_), .B1(KEYINPUT111), .B2(KEYINPUT52), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n814_), .A2(new_n817_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n812_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT53), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n812_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1339gat));
  INV_X1    g622(.A(new_n493_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n490_), .A2(new_n492_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n765_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n500_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n584_), .B2(new_n579_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT115), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n829_), .C1(new_n584_), .C2(new_n579_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n501_), .A2(new_n581_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n570_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n607_), .A2(new_n561_), .B1(new_n835_), .B2(new_n577_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n573_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n563_), .A2(new_n571_), .A3(KEYINPUT55), .A4(new_n565_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n590_), .A2(new_n576_), .A3(new_n534_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT12), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n552_), .A2(new_n562_), .B1(new_n841_), .B2(new_n568_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT55), .B1(new_n842_), .B2(new_n565_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n509_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT56), .B(new_n509_), .C1(new_n839_), .C2(new_n843_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n834_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n831_), .B(new_n833_), .C1(new_n848_), .C2(KEYINPUT114), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n766_), .A2(new_n584_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n847_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n572_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n854_), .B2(new_n509_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n850_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n629_), .B1(new_n849_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n581_), .B(new_n829_), .C1(new_n851_), .C2(new_n855_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT116), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n632_), .B1(new_n862_), .B2(KEYINPUT58), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(KEYINPUT116), .A3(new_n864_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n859_), .A2(new_n860_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n831_), .A2(new_n833_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n848_), .A2(KEYINPUT114), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n860_), .B(new_n666_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n646_), .B1(new_n866_), .B2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n632_), .A2(new_n766_), .A3(new_n586_), .A4(new_n646_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT54), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT113), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n876_), .A3(KEYINPUT54), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n587_), .B(new_n696_), .C1(new_n631_), .C2(new_n630_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .A4(new_n766_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT112), .B1(new_n873_), .B2(KEYINPUT54), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n875_), .A2(new_n877_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n872_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n655_), .A2(new_n656_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n259_), .A3(new_n658_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G113gat), .B1(new_n887_), .B2(new_n501_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n829_), .A2(new_n581_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n711_), .A2(new_n865_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n666_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(KEYINPUT57), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n696_), .B1(new_n896_), .B2(new_n870_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(KEYINPUT119), .B(new_n696_), .C1(new_n896_), .C2(new_n870_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n883_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n886_), .A2(KEYINPUT118), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n886_), .A2(KEYINPUT118), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI22_X1  g705(.A1(new_n887_), .A2(new_n889_), .B1(new_n901_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n766_), .A2(KEYINPUT120), .ZN(new_n909_));
  MUX2_X1   g708(.A(KEYINPUT120), .B(new_n909_), .S(G113gat), .Z(new_n910_));
  AOI21_X1  g709(.A(new_n888_), .B1(new_n908_), .B2(new_n910_), .ZN(G1340gat));
  OAI21_X1  g710(.A(G120gat), .B1(new_n907_), .B2(new_n586_), .ZN(new_n912_));
  INV_X1    g711(.A(G120gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n887_), .B(new_n914_), .C1(KEYINPUT60), .C2(new_n913_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(G1341gat));
  OAI21_X1  g715(.A(G127gat), .B1(new_n907_), .B2(new_n696_), .ZN(new_n917_));
  INV_X1    g716(.A(G127gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n887_), .A2(new_n918_), .A3(new_n646_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1342gat));
  OAI21_X1  g719(.A(G134gat), .B1(new_n907_), .B2(new_n632_), .ZN(new_n921_));
  INV_X1    g720(.A(G134gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n887_), .A2(new_n922_), .A3(new_n666_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1343gat));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925_));
  NOR4_X1   g724(.A1(new_n658_), .A2(new_n437_), .A3(new_n654_), .A4(new_n450_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n925_), .B1(new_n884_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n875_), .A2(new_n877_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n881_), .A2(new_n882_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n897_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(KEYINPUT121), .A3(new_n926_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n766_), .B1(new_n928_), .B2(new_n933_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT122), .B(G141gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1344gat));
  AOI21_X1  g735(.A(new_n586_), .B1(new_n928_), .B2(new_n933_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT123), .B(G148gat), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n937_), .B(new_n939_), .ZN(G1345gat));
  AOI21_X1  g739(.A(new_n696_), .B1(new_n928_), .B2(new_n933_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT61), .B(G155gat), .Z(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT124), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(KEYINPUT125), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n941_), .B(new_n944_), .ZN(G1346gat));
  NAND2_X1  g744(.A1(new_n928_), .A2(new_n933_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n946_), .A2(new_n216_), .A3(new_n666_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n632_), .B1(new_n928_), .B2(new_n933_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n216_), .B2(new_n948_), .ZN(G1347gat));
  NAND2_X1  g748(.A1(new_n330_), .A2(new_n654_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n449_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n899_), .A2(new_n900_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n931_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  OAI211_X1 g754(.A(KEYINPUT62), .B(G169gat), .C1(new_n955_), .C2(new_n766_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n901_), .A2(new_n766_), .A3(new_n952_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n286_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n958_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n956_), .A2(new_n959_), .A3(new_n960_), .ZN(G1348gat));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962_));
  AOI21_X1  g761(.A(G176gat), .B1(new_n954_), .B2(new_n587_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n884_), .A2(new_n449_), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n950_), .A2(new_n298_), .A3(new_n586_), .ZN(new_n965_));
  AND2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n962_), .B1(new_n963_), .B2(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n964_), .A2(new_n965_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n901_), .A2(new_n586_), .A3(new_n952_), .ZN(new_n969_));
  OAI211_X1 g768(.A(KEYINPUT126), .B(new_n968_), .C1(new_n969_), .C2(G176gat), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n967_), .A2(new_n970_), .ZN(G1349gat));
  NOR2_X1   g770(.A1(new_n950_), .A2(new_n696_), .ZN(new_n972_));
  AOI21_X1  g771(.A(G183gat), .B1(new_n964_), .B2(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n696_), .A2(new_n340_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n954_), .B2(new_n974_), .ZN(G1350gat));
  OAI21_X1  g774(.A(G190gat), .B1(new_n955_), .B2(new_n632_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n954_), .A2(new_n339_), .A3(new_n666_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1351gat));
  NOR4_X1   g777(.A1(new_n658_), .A2(new_n437_), .A3(new_n414_), .A4(new_n259_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n932_), .A2(new_n979_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(new_n766_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(new_n364_), .ZN(G1352gat));
  NOR2_X1   g781(.A1(new_n980_), .A2(new_n586_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(new_n366_), .ZN(G1353gat));
  NOR2_X1   g783(.A1(new_n980_), .A2(new_n696_), .ZN(new_n985_));
  NOR3_X1   g784(.A1(new_n985_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986_));
  XOR2_X1   g785(.A(KEYINPUT63), .B(G211gat), .Z(new_n987_));
  AOI21_X1  g786(.A(new_n986_), .B1(new_n985_), .B2(new_n987_), .ZN(G1354gat));
  OAI21_X1  g787(.A(G218gat), .B1(new_n980_), .B2(new_n632_), .ZN(new_n989_));
  OR2_X1    g788(.A1(new_n629_), .A2(G218gat), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n980_), .B2(new_n990_), .ZN(G1355gat));
endmodule


