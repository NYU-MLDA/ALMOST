//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT88), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT89), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT89), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n212_), .A3(new_n209_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n205_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n204_), .B(KEYINPUT1), .Z(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(new_n203_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n208_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G127gat), .B(G134gat), .Z(new_n223_));
  XOR2_X1   g022(.A(G113gat), .B(G120gat), .Z(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(KEYINPUT98), .B(new_n225_), .C1(new_n214_), .C2(new_n221_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n214_), .A2(new_n221_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n230_), .A2(KEYINPUT98), .A3(new_n231_), .A4(new_n225_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n225_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n237_), .B2(new_n227_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G1gat), .B(G29gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G85gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n236_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n234_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n238_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G8gat), .B(G36gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT18), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G64gat), .B(G92gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT83), .B(G183gat), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT25), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263_));
  INV_X1    g062(.A(G190gat), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n263_), .A2(G183gat), .B1(new_n264_), .B2(KEYINPUT26), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n257_), .A2(new_n259_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT23), .ZN(new_n268_));
  INV_X1    g067(.A(G169gat), .ZN(new_n269_));
  INV_X1    g068(.A(G176gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT24), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(KEYINPUT24), .A3(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n266_), .A2(new_n268_), .A3(new_n272_), .A4(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n256_), .A2(new_n264_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n268_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT22), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT85), .B1(new_n278_), .B2(G169gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT86), .B(G176gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT22), .B(G169gat), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n279_), .B(new_n280_), .C1(new_n281_), .C2(KEYINPUT85), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n273_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G204gat), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G197gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT21), .ZN(new_n290_));
  XOR2_X1   g089(.A(G211gat), .B(G218gat), .Z(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n289_), .A2(KEYINPUT93), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT93), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT21), .B1(new_n286_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(KEYINPUT21), .A3(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n284_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n264_), .A2(KEYINPUT26), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n260_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n268_), .B1(new_n271_), .B2(new_n306_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n268_), .B1(G183gat), .B2(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n281_), .A2(new_n280_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n273_), .A3(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n310_), .A2(new_n296_), .A3(new_n297_), .A4(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n299_), .A2(KEYINPUT20), .A3(new_n302_), .A4(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n309_), .B2(new_n308_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n298_), .B2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n275_), .A2(new_n296_), .A3(new_n297_), .A4(new_n283_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n302_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n255_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n254_), .A3(new_n315_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT96), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT27), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT96), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n323_), .A2(new_n327_), .A3(new_n254_), .A4(new_n315_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n319_), .A2(new_n302_), .A3(new_n320_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT102), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT102), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n319_), .A2(new_n332_), .A3(new_n320_), .A4(new_n302_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n299_), .A2(KEYINPUT20), .A3(new_n314_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n331_), .B(new_n333_), .C1(new_n302_), .C2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n255_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT27), .A3(new_n324_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n250_), .A2(new_n329_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G43gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n284_), .B(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n341_), .A2(new_n226_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n226_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(G15gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT31), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n342_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n298_), .B1(new_n222_), .B2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(G233gat), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G78gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G106gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n355_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  XOR2_X1   g162(.A(G22gat), .B(G50gat), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT91), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n222_), .A2(new_n354_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n222_), .B2(new_n354_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n365_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n362_), .A2(new_n363_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n363_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n362_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n363_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n353_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n352_), .B(new_n375_), .C1(new_n379_), .C2(new_n378_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n338_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n323_), .A2(new_n315_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n335_), .A2(KEYINPUT103), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT103), .B1(new_n335_), .B2(new_n385_), .ZN(new_n387_));
  OAI221_X1 g186(.A(new_n249_), .B1(new_n384_), .B2(new_n385_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n325_), .A2(new_n328_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT97), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n229_), .A2(new_n234_), .A3(new_n232_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n237_), .A2(new_n235_), .A3(new_n227_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n244_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT101), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT101), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n392_), .A2(new_n396_), .A3(new_n244_), .A4(new_n393_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n248_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n325_), .A2(KEYINPUT97), .A3(new_n328_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n391_), .A2(new_n398_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n248_), .A2(new_n399_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT100), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n388_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n380_), .A2(new_n352_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n383_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G1gat), .B(G8gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G22gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n345_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G15gat), .A2(G22gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G1gat), .A2(G8gat), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n413_), .A2(new_n414_), .B1(KEYINPUT14), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n411_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G29gat), .B(G36gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(KEYINPUT76), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(KEYINPUT76), .ZN(new_n421_));
  XOR2_X1   g220(.A(G43gat), .B(G50gat), .Z(new_n422_));
  OR3_X1    g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT15), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT15), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n417_), .A2(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G229gat), .A2(G233gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n430_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n417_), .A2(new_n425_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G113gat), .B(G141gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G169gat), .B(G197gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n432_), .A2(new_n436_), .A3(KEYINPUT82), .A4(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n436_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n439_), .B(KEYINPUT81), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G64gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G57gat), .ZN(new_n451_));
  INV_X1    g250(.A(G57gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT68), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT68), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G71gat), .B(G78gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n463_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT68), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT68), .B1(new_n451_), .B2(new_n453_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT11), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT69), .B1(new_n470_), .B2(new_n461_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n465_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT71), .B1(new_n467_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT9), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT65), .B(G92gat), .Z(new_n477_));
  INV_X1    g276(.A(G85gat), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n475_), .B(new_n476_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n478_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT66), .B1(new_n482_), .B2(KEYINPUT9), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  AND2_X1   g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(KEYINPUT9), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT6), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n488_), .A2(new_n489_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n487_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496_));
  INV_X1    g295(.A(G99gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n489_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n491_), .A2(new_n493_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n496_), .A2(new_n497_), .A3(new_n489_), .A4(KEYINPUT67), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n485_), .A2(new_n484_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n506_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT8), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT70), .B1(new_n513_), .B2(new_n507_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n495_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n466_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n471_), .A2(new_n472_), .A3(new_n465_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n474_), .A2(new_n515_), .A3(KEYINPUT12), .A4(new_n519_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n513_), .A2(new_n507_), .B1(new_n487_), .B2(new_n494_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n516_), .A2(new_n521_), .A3(new_n517_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT64), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n520_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G120gat), .B(G148gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT73), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT74), .Z(new_n539_));
  AND3_X1   g338(.A1(new_n530_), .A2(new_n533_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n546_), .B(new_n547_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(G231gat), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n516_), .A2(new_n517_), .A3(new_n417_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n417_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n552_));
  INV_X1    g351(.A(G233gat), .ZN(new_n553_));
  OR4_X1    g352(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n551_), .A2(new_n552_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT17), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n518_), .A3(KEYINPUT17), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT80), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .A4(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT36), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n515_), .A2(new_n428_), .A3(new_n427_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n521_), .A2(new_n425_), .B1(new_n580_), .B2(new_n579_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n575_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n572_), .A2(new_n573_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n590_), .A3(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT37), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n567_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR4_X1   g396(.A1(new_n408_), .A2(new_n449_), .A3(new_n549_), .A4(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n249_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n592_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n408_), .A2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n549_), .A2(new_n449_), .A3(new_n567_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n250_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n601_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n607_), .A3(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(G8gat), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n329_), .A2(new_n337_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n598_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n606_), .B2(new_n611_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n613_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g417(.A(new_n606_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n353_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G15gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT104), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n623_), .A3(G15gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(KEYINPUT41), .A3(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n598_), .A2(new_n345_), .A3(new_n353_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(new_n622_), .B2(new_n624_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(new_n380_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n598_), .A2(new_n412_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G22gat), .B1(new_n606_), .B2(new_n380_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT42), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT42), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT105), .ZN(G1327gat));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n593_), .A2(new_n595_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT107), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n408_), .B2(new_n638_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n638_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n403_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n401_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT97), .B1(new_n325_), .B2(new_n328_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n400_), .A2(new_n398_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n406_), .B1(new_n650_), .B2(new_n388_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n643_), .B(new_n640_), .C1(new_n651_), .C2(new_n383_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n642_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n567_), .ZN(new_n654_));
  OR4_X1    g453(.A1(KEYINPUT106), .A2(new_n549_), .A3(new_n449_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n549_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n448_), .A3(new_n567_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT106), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n653_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n642_), .A2(new_n652_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT108), .B1(new_n663_), .B2(KEYINPUT44), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n665_), .A3(new_n661_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n637_), .B1(new_n667_), .B2(new_n249_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n405_), .A2(new_n407_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n383_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n654_), .A2(new_n592_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(new_n448_), .A3(new_n656_), .A4(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(G29gat), .A3(new_n250_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT109), .B1(new_n668_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n676_));
  INV_X1    g475(.A(new_n674_), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n250_), .B(new_n662_), .C1(new_n664_), .C2(new_n666_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n676_), .B(new_n677_), .C1(new_n678_), .C2(new_n637_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n663_), .A2(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n665_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n663_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n612_), .B(new_n685_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G36gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n673_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n611_), .A2(G36gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n692_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT45), .B1(new_n673_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n681_), .A2(new_n682_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n684_), .B1(new_n689_), .B2(new_n699_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n683_), .B(new_n698_), .C1(new_n688_), .C2(G36gat), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  AOI21_X1  g501(.A(G43gat), .B1(new_n690_), .B2(new_n353_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n353_), .A2(G43gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n667_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1330gat));
  AOI21_X1  g506(.A(G50gat), .B1(new_n690_), .B2(new_n630_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n630_), .A2(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n667_), .B2(new_n709_), .ZN(G1331gat));
  NOR4_X1   g509(.A1(new_n408_), .A2(new_n448_), .A3(new_n656_), .A4(new_n597_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n452_), .A3(new_n249_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n656_), .A2(new_n448_), .A3(new_n567_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n604_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(new_n249_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n712_), .B1(new_n715_), .B2(new_n452_), .ZN(G1332gat));
  AOI21_X1  g515(.A(new_n450_), .B1(new_n714_), .B2(new_n612_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT48), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n711_), .A2(new_n450_), .A3(new_n612_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1333gat));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n711_), .A2(new_n721_), .A3(new_n353_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n714_), .A2(new_n353_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(G71gat), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT112), .Z(G1334gat));
  AOI21_X1  g527(.A(new_n359_), .B1(new_n714_), .B2(new_n630_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n380_), .A2(G78gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT114), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n711_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1335gat));
  AND4_X1   g534(.A1(new_n671_), .A2(new_n449_), .A3(new_n549_), .A4(new_n672_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n478_), .A3(new_n249_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n549_), .A2(new_n449_), .A3(new_n567_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n642_), .B2(new_n652_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(new_n249_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n740_), .B2(new_n478_), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n736_), .B2(new_n612_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n611_), .A2(new_n477_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n739_), .B2(new_n743_), .ZN(G1337gat));
  NAND2_X1  g543(.A1(new_n353_), .A2(new_n488_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT115), .B1(new_n736_), .B2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n739_), .A2(new_n353_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n497_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g549(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n739_), .A2(new_n630_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G106gat), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n736_), .A2(new_n489_), .A3(new_n630_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n751_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n751_), .ZN(new_n760_));
  AOI211_X1 g559(.A(new_n757_), .B(new_n760_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  NAND4_X1  g561(.A1(new_n596_), .A2(new_n449_), .A3(new_n545_), .A4(new_n548_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n530_), .A2(new_n533_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(new_n537_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n448_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n520_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n532_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n530_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n520_), .A2(new_n525_), .A3(new_n529_), .A4(KEYINPUT55), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n537_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n768_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n439_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(KEYINPUT117), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n781_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n434_), .A2(new_n431_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n783_), .A2(new_n784_), .B1(new_n429_), .B2(new_n785_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n782_), .A2(new_n786_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n542_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n592_), .B1(new_n779_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n767_), .A2(new_n448_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n537_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n788_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n767_), .A2(new_n787_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n799_), .B(KEYINPUT58), .C1(new_n794_), .C2(new_n795_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n643_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n792_), .A2(new_n798_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n765_), .B1(new_n805_), .B2(new_n567_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n612_), .A2(new_n250_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n381_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n448_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n802_), .A2(new_n643_), .A3(new_n803_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n797_), .B2(new_n592_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT118), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n792_), .A2(new_n815_), .A3(new_n804_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n798_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n765_), .B1(new_n817_), .B2(new_n567_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n806_), .B2(new_n809_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n448_), .A2(G113gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n811_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(new_n820_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n549_), .B(new_n822_), .C1(new_n818_), .C2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G120gat), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n830_));
  AOI21_X1  g629(.A(G120gat), .B1(new_n549_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(G120gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(KEYINPUT120), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(KEYINPUT120), .B2(new_n831_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n810_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n829_), .A2(new_n838_), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1341gat));
  NAND3_X1  g639(.A1(new_n821_), .A2(new_n654_), .A3(new_n822_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G127gat), .ZN(new_n842_));
  INV_X1    g641(.A(new_n810_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n567_), .A2(G127gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(G1342gat));
  NAND3_X1  g644(.A1(new_n821_), .A2(new_n643_), .A3(new_n822_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G134gat), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n592_), .A2(G134gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n843_), .B2(new_n848_), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n806_), .A2(new_n382_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n807_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n449_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n656_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g654(.A1(new_n851_), .A2(new_n567_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT61), .B(G155gat), .Z(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  INV_X1    g657(.A(G162gat), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n851_), .A2(new_n859_), .A3(new_n638_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n851_), .B2(new_n592_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n861_), .A2(KEYINPUT122), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(KEYINPUT122), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(G1347gat));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n269_), .B1(new_n865_), .B2(KEYINPUT62), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n611_), .A2(new_n249_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n353_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n630_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n819_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n870_), .B2(new_n449_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI221_X1 g672(.A(new_n866_), .B1(new_n865_), .B2(KEYINPUT62), .C1(new_n870_), .C2(new_n449_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n870_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n281_), .A3(new_n448_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n874_), .A3(new_n876_), .ZN(G1348gat));
  INV_X1    g676(.A(new_n806_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n380_), .ZN(new_n879_));
  NOR4_X1   g678(.A1(new_n879_), .A2(new_n270_), .A3(new_n656_), .A4(new_n868_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n549_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n280_), .ZN(G1349gat));
  NOR3_X1   g681(.A1(new_n870_), .A2(new_n303_), .A3(new_n567_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n868_), .A2(new_n567_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n878_), .A2(new_n380_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT124), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n883_), .B1(new_n256_), .B2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n870_), .B2(new_n638_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n603_), .A2(new_n260_), .A3(new_n304_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n870_), .B2(new_n889_), .ZN(G1351gat));
  NAND2_X1  g689(.A1(new_n850_), .A2(new_n867_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n449_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n285_), .ZN(G1352gat));
  INV_X1    g692(.A(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n549_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT125), .B(G204gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1353gat));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n567_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n891_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(G211gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n850_), .A2(new_n903_), .A3(new_n867_), .A4(new_n899_), .ZN(new_n904_));
  AND4_X1   g703(.A1(new_n898_), .A2(new_n901_), .A3(new_n902_), .A4(new_n904_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n901_), .A2(new_n904_), .B1(new_n898_), .B2(new_n902_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1354gat));
  XNOR2_X1  g706(.A(KEYINPUT127), .B(G218gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n891_), .A2(new_n638_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n894_), .A2(new_n603_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(G1355gat));
endmodule


