//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(new_n205_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  OAI221_X1 g013(.A(new_n212_), .B1(G85gat), .B2(G92gat), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(G106gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n211_), .A2(new_n218_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n207_), .A2(new_n221_), .A3(new_n210_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT66), .B1(new_n223_), .B2(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G85gat), .B(G92gat), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(new_n232_), .B2(new_n208_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT68), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(new_n231_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(new_n206_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n236_), .B(KEYINPUT8), .C1(new_n239_), .C2(new_n227_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n211_), .A2(new_n232_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n241_), .A2(KEYINPUT72), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT72), .B1(new_n241_), .B2(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n226_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G29gat), .B(G36gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G43gat), .B(G50gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT15), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n241_), .A2(new_n244_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n226_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(KEYINPUT75), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT35), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n252_), .A2(new_n254_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n255_), .B(new_n260_), .C1(new_n261_), .C2(KEYINPUT35), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT36), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G190gat), .B(G218gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT76), .ZN(new_n265_));
  XOR2_X1   g064(.A(G134gat), .B(G162gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n252_), .A2(KEYINPUT75), .A3(new_n254_), .A4(new_n259_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n262_), .A2(new_n263_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n255_), .A2(new_n260_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT35), .B1(new_n252_), .B2(new_n254_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n267_), .B(KEYINPUT36), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(new_n274_), .A3(KEYINPUT37), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n273_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n272_), .B2(KEYINPUT77), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT77), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n262_), .A2(new_n279_), .A3(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n269_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT37), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n276_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G8gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT78), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT78), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  INV_X1    g088(.A(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT14), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n286_), .A2(new_n292_), .A3(new_n289_), .A4(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G231gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT69), .B(G71gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(G78gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(G78gat), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n304_), .B(new_n305_), .C1(KEYINPUT11), .C2(new_n299_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n302_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n298_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G127gat), .B(G155gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G183gat), .B(G211gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT17), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(KEYINPUT17), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n308_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n308_), .A2(new_n315_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n284_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT80), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n247_), .A2(KEYINPUT12), .A3(new_n307_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n235_), .A2(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n324_), .A2(new_n307_), .A3(new_n225_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT12), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n307_), .B1(new_n324_), .B2(new_n225_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n302_), .B(new_n306_), .Z(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n226_), .A3(new_n253_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(new_n327_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n330_), .B1(new_n333_), .B2(new_n323_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n323_), .B1(new_n332_), .B2(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT71), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G120gat), .B(G148gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT5), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n329_), .A2(new_n334_), .A3(new_n336_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT73), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n335_), .B(new_n330_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n329_), .A4(new_n341_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n329_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n340_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(KEYINPUT13), .A3(new_n349_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n296_), .A2(new_n250_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT81), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n296_), .A2(new_n250_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G229gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n296_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n356_), .B1(new_n362_), .B2(new_n251_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G141gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G169gat), .B(G197gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  OR2_X1    g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n354_), .A2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(KEYINPUT88), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT85), .B(G197gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(G204gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(G211gat), .B(G218gat), .Z(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(KEYINPUT21), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT87), .B1(new_n376_), .B2(KEYINPUT21), .ZN(new_n380_));
  AND2_X1   g179(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(G204gat), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n374_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT21), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G204gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n390_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT86), .B1(new_n390_), .B2(G197gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n377_), .B1(new_n394_), .B2(KEYINPUT21), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n379_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n372_), .A2(KEYINPUT88), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398_));
  INV_X1    g197(.A(G141gat), .ZN(new_n399_));
  INV_X1    g198(.A(G148gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n401_), .A2(new_n403_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G155gat), .B(G162gat), .Z(new_n407_));
  INV_X1    g206(.A(G155gat), .ZN(new_n408_));
  INV_X1    g207(.A(G162gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT1), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT1), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G155gat), .A3(G162gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n409_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G141gat), .B(G148gat), .Z(new_n415_));
  AOI22_X1  g214(.A1(new_n406_), .A2(new_n407_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n397_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n373_), .B1(new_n396_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n386_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n420_));
  AOI211_X1 g219(.A(KEYINPUT87), .B(KEYINPUT21), .C1(new_n383_), .C2(new_n384_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n395_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n378_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n418_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n373_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n419_), .B2(new_n426_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n419_), .A2(new_n426_), .A3(KEYINPUT89), .A4(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n406_), .A2(new_n407_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n414_), .A2(new_n415_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n417_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT28), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n416_), .A2(new_n438_), .A3(new_n417_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G22gat), .B(G50gat), .Z(new_n440_));
  AND3_X1   g239(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n433_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n419_), .A2(new_n426_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n427_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n443_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n419_), .A2(new_n426_), .A3(KEYINPUT90), .A4(new_n427_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n428_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n444_), .A2(new_n445_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n443_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT91), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G226gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT19), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT82), .B(G190gat), .ZN(new_n462_));
  INV_X1    g261(.A(G183gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G183gat), .A2(G190gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT23), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n468_));
  AOI21_X1  g267(.A(G176gat), .B1(new_n468_), .B2(KEYINPUT22), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(G169gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT25), .B(G183gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT26), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G190gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n462_), .B2(KEYINPUT26), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n462_), .A2(new_n476_), .A3(KEYINPUT26), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n465_), .B(KEYINPUT23), .Z(new_n481_));
  NOR2_X1   g280(.A1(G169gat), .A2(G176gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G169gat), .ZN(new_n485_));
  INV_X1    g284(.A(G176gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT24), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n484_), .B1(new_n487_), .B2(new_n482_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n471_), .B1(new_n480_), .B2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(KEYINPUT92), .B(KEYINPUT20), .C1(new_n423_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n481_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(G183gat), .B2(G190gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n485_), .A2(new_n486_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT22), .B(G169gat), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n486_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT26), .B(G190gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n481_), .B1(new_n472_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n488_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n494_), .A2(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n423_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n462_), .A2(new_n476_), .A3(KEYINPUT26), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n472_), .B(new_n474_), .C1(new_n505_), .C2(new_n477_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n506_), .A2(new_n489_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n396_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT92), .B1(new_n508_), .B2(KEYINPUT20), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n461_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G8gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT18), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT93), .B1(new_n396_), .B2(new_n507_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n423_), .A2(new_n517_), .A3(new_n491_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n461_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n396_), .B2(new_n501_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n510_), .A2(new_n515_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT27), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n522_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n461_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n521_), .B1(new_n396_), .B2(new_n507_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(KEYINPUT92), .B1(new_n423_), .B2(new_n502_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n508_), .A2(KEYINPUT20), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n532_), .A3(new_n520_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n515_), .B1(new_n527_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n525_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n520_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n514_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT27), .B1(new_n538_), .B2(new_n524_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n459_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n434_), .A2(new_n435_), .ZN(new_n542_));
  INV_X1    g341(.A(G134gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(G127gat), .ZN(new_n544_));
  INV_X1    g343(.A(G127gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G134gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G120gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G113gat), .ZN(new_n549_));
  INV_X1    g348(.A(G113gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G120gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n544_), .A2(new_n546_), .A3(new_n549_), .A4(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n542_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT95), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(KEYINPUT4), .A3(new_n559_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT94), .ZN(new_n563_));
  INV_X1    g362(.A(new_n558_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n557_), .A2(new_n559_), .A3(new_n565_), .A4(KEYINPUT4), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n557_), .A2(KEYINPUT4), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G29gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G85gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT0), .B(G57gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  AND3_X1   g371(.A1(new_n561_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n561_), .B2(new_n568_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT99), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n561_), .A2(new_n568_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n561_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G71gat), .B(G99gat), .ZN(new_n584_));
  INV_X1    g383(.A(G43gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n507_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n555_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G227gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(G15gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT30), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT31), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n588_), .B(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n583_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n541_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n445_), .B1(new_n444_), .B2(new_n452_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT91), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n583_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n524_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n515_), .B1(new_n510_), .B2(new_n523_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI22_X1  g402(.A1(new_n603_), .A2(KEYINPUT27), .B1(new_n534_), .B2(new_n525_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n597_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n582_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n540_), .A3(KEYINPUT100), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n527_), .A2(new_n533_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n515_), .A2(KEYINPUT32), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n608_), .A2(new_n609_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(KEYINPUT98), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n510_), .A3(new_n523_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n580_), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT97), .B1(new_n557_), .B2(new_n559_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n558_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n557_), .A2(KEYINPUT97), .A3(new_n559_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n572_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n563_), .A2(new_n558_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n616_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n580_), .A2(new_n615_), .A3(new_n614_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n623_), .A2(new_n524_), .A3(new_n538_), .A4(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n613_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n459_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n605_), .A2(new_n607_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n594_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n596_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n371_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n321_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(KEYINPUT38), .A3(new_n290_), .A4(new_n582_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n267_), .A2(new_n263_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n272_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n630_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n637_), .A2(new_n319_), .A3(new_n370_), .A4(new_n354_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n638_), .B2(new_n583_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n321_), .A2(new_n631_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n582_), .A2(new_n290_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n633_), .A2(new_n639_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n638_), .A2(new_n540_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(new_n291_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT102), .B(G8gat), .C1(new_n638_), .C2(new_n540_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(KEYINPUT39), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n647_), .B(new_n652_), .C1(new_n648_), .C2(new_n291_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n632_), .A2(new_n291_), .A3(new_n604_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n651_), .A2(KEYINPUT40), .A3(new_n653_), .A4(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1325gat));
  NAND3_X1  g458(.A1(new_n632_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT103), .ZN(new_n661_));
  OAI21_X1  g460(.A(G15gat), .B1(new_n638_), .B2(new_n629_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n663_), .A3(new_n664_), .ZN(G1326gat));
  OAI21_X1  g464(.A(G22gat), .B1(new_n638_), .B2(new_n459_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n641_), .A2(G22gat), .A3(new_n459_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT104), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n671_), .A3(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n282_), .A2(new_n319_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n371_), .A2(new_n630_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n582_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n630_), .B2(new_n284_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n275_), .B1(new_n636_), .B2(KEYINPUT37), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n606_), .A2(new_n540_), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n682_), .A2(new_n597_), .B1(new_n459_), .B2(new_n626_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n594_), .B1(new_n683_), .B2(new_n607_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n680_), .B(new_n681_), .C1(new_n684_), .C2(new_n596_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n319_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n354_), .A2(new_n687_), .A3(new_n370_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AND4_X1   g488(.A1(KEYINPUT106), .A2(new_n686_), .A3(KEYINPUT44), .A4(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n679_), .B2(new_n685_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT106), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  INV_X1    g493(.A(new_n678_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n596_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n606_), .A2(new_n540_), .A3(KEYINPUT100), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT100), .B1(new_n606_), .B2(new_n540_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n458_), .B1(new_n613_), .B2(new_n625_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n700_), .B2(new_n594_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n695_), .B1(new_n701_), .B2(new_n681_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n630_), .A2(KEYINPUT43), .A3(new_n284_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n689_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n693_), .B1(new_n694_), .B2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n582_), .A2(G29gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n677_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  XNOR2_X1  g506(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n540_), .B1(new_n704_), .B2(new_n694_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n631_), .A2(new_n674_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n540_), .A2(G36gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT45), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n676_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n708_), .B1(new_n711_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n708_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n718_), .B(new_n721_), .C1(new_n710_), .C2(G36gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1329gat));
  NOR2_X1   g522(.A1(new_n629_), .A2(new_n585_), .ZN(new_n724_));
  OAI221_X1 g523(.A(new_n724_), .B1(KEYINPUT44), .B2(new_n691_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n585_), .B1(new_n712_), .B2(new_n629_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT47), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n729_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n676_), .B2(new_n458_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n458_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n705_), .B2(new_n733_), .ZN(G1331gat));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n582_), .B2(KEYINPUT110), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n352_), .A2(new_n353_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n370_), .A2(new_n687_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n637_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n736_), .B(new_n739_), .C1(KEYINPUT110), .C2(new_n735_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n321_), .A2(new_n737_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT108), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n630_), .A2(new_n370_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(KEYINPUT109), .ZN(new_n744_));
  INV_X1    g543(.A(new_n370_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n701_), .A2(KEYINPUT109), .A3(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n582_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n740_), .B1(new_n748_), .B2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g548(.A(G64gat), .B1(new_n739_), .B2(new_n540_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT48), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n742_), .A2(new_n747_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n540_), .A2(G64gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n739_), .B2(new_n629_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT49), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n629_), .A2(G71gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n752_), .B2(new_n757_), .ZN(G1334gat));
  OAI21_X1  g557(.A(G78gat), .B1(new_n739_), .B2(new_n459_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n459_), .A2(G78gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n752_), .B2(new_n762_), .ZN(G1335gat));
  NAND3_X1  g562(.A1(new_n737_), .A2(new_n687_), .A3(new_n745_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n686_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n583_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n675_), .A2(new_n354_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n747_), .A2(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n583_), .A2(G85gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n766_), .B2(new_n540_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n540_), .A2(G92gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n769_), .B2(new_n773_), .ZN(G1337gat));
  NOR2_X1   g573(.A1(new_n629_), .A2(new_n220_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n768_), .B(new_n775_), .C1(new_n744_), .C2(new_n746_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n686_), .A2(new_n594_), .A3(new_n765_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G99gat), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(G1338gat));
  AOI211_X1 g585(.A(new_n459_), .B(new_n764_), .C1(new_n679_), .C2(new_n685_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT114), .B1(new_n787_), .B2(new_n229_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n686_), .A2(new_n458_), .A3(new_n765_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(KEYINPUT52), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n459_), .A2(G106gat), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n788_), .A2(KEYINPUT52), .B1(new_n769_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n793_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n769_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n798_), .A2(new_n794_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n792_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n803_), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n358_), .A2(new_n360_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n367_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n806_), .A2(new_n807_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT117), .B1(new_n805_), .B2(new_n367_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n808_), .A2(new_n809_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n350_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n323_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n329_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n322_), .A2(new_n328_), .A3(KEYINPUT55), .A4(new_n323_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n340_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n818_), .B2(KEYINPUT116), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n341_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT115), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n347_), .B(new_n370_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n811_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n282_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n282_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n823_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n282_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n810_), .A2(new_n347_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n820_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n832_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n831_), .A2(KEYINPUT58), .A3(new_n833_), .A4(new_n834_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n681_), .A3(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n826_), .A2(new_n829_), .A3(new_n830_), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n687_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n284_), .A2(new_n354_), .A3(new_n842_), .A4(new_n738_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n352_), .A2(new_n353_), .A3(new_n738_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT54), .B1(new_n844_), .B2(new_n681_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n846_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n541_), .A2(new_n583_), .A3(new_n629_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(KEYINPUT119), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  INV_X1    g649(.A(new_n846_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n840_), .B2(new_n687_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n848_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n850_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n849_), .A2(new_n854_), .A3(new_n550_), .A4(new_n370_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(KEYINPUT59), .A3(new_n848_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n745_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n859_), .B2(new_n550_), .ZN(G1340gat));
  AOI21_X1  g659(.A(new_n354_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT120), .B(G120gat), .Z(new_n862_));
  NAND2_X1  g661(.A1(new_n849_), .A2(new_n854_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n354_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(KEYINPUT60), .B2(new_n862_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n861_), .A2(new_n862_), .B1(new_n863_), .B2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g665(.A(new_n687_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n319_), .A2(new_n545_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n867_), .A2(new_n545_), .B1(new_n863_), .B2(new_n868_), .ZN(G1342gat));
  AOI21_X1  g668(.A(new_n284_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n636_), .A2(new_n543_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n870_), .A2(new_n543_), .B1(new_n863_), .B2(new_n871_), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n459_), .A2(new_n594_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n604_), .A3(new_n583_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n370_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n737_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT121), .B(G148gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1345gat));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n847_), .A2(new_n319_), .A3(new_n875_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n877_), .A2(KEYINPUT122), .A3(new_n319_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT122), .B1(new_n877_), .B2(new_n319_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n852_), .A2(new_n885_), .A3(new_n687_), .A4(new_n876_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n883_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1346gat));
  INV_X1    g692(.A(new_n877_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G162gat), .B1(new_n894_), .B2(new_n284_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n877_), .A2(new_n409_), .A3(new_n636_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n595_), .A2(new_n540_), .A3(new_n458_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n847_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n745_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n901_), .B2(new_n485_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n496_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT62), .B(G169gat), .C1(new_n900_), .C2(new_n745_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n900_), .A2(new_n354_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n486_), .ZN(G1349gat));
  NOR3_X1   g706(.A1(new_n900_), .A2(new_n687_), .A3(new_n472_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n900_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n319_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n463_), .B2(new_n910_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n900_), .B2(new_n284_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n636_), .A2(new_n498_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n900_), .B2(new_n913_), .ZN(G1351gat));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n874_), .A2(new_n540_), .A3(new_n582_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n847_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n916_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT123), .B1(new_n852_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G197gat), .B1(new_n920_), .B2(new_n370_), .ZN(new_n921_));
  INV_X1    g720(.A(G197gat), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n922_), .B(new_n745_), .C1(new_n917_), .C2(new_n919_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1352gat));
  AOI21_X1  g723(.A(new_n915_), .B1(new_n847_), .B2(new_n916_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n852_), .A2(KEYINPUT123), .A3(new_n918_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n737_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n390_), .A2(KEYINPUT124), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT125), .Z(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n920_), .A2(new_n737_), .A3(new_n929_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1353gat));
  NOR3_X1   g732(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n934_));
  AOI211_X1 g733(.A(new_n934_), .B(new_n687_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n920_), .A2(new_n937_), .A3(new_n935_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1354gat));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n920_), .A2(new_n942_), .A3(new_n636_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n284_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n942_), .B2(new_n944_), .ZN(G1355gat));
endmodule


