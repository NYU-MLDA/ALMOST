//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(KEYINPUT80), .B(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  OR2_X1    g002(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(G190gat), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT79), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT79), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G183gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT25), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n203_), .B(new_n206_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(new_n214_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n221_), .A2(KEYINPUT24), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n213_), .A2(new_n218_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT82), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT23), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n214_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n214_), .A2(new_n235_), .A3(KEYINPUT23), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n208_), .A2(new_n210_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(new_n202_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n229_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n226_), .A2(new_n227_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n227_), .B1(new_n226_), .B2(new_n241_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT31), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT31), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT30), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G15gat), .B(G43gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT85), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(G227gat), .A3(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(G227gat), .ZN(new_n262_));
  INV_X1    g061(.A(G233gat), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n257_), .B(new_n259_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G71gat), .B(G99gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n266_), .A3(new_n264_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n252_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(new_n252_), .A3(new_n269_), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n249_), .A2(new_n250_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n250_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n270_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n248_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT95), .B(G78gat), .ZN(new_n277_));
  INV_X1    g076(.A(G106gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G197gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G197gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n284_), .A3(KEYINPUT91), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n285_), .B(KEYINPUT21), .C1(KEYINPUT91), .C2(new_n282_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n288_), .A2(new_n282_), .A3(new_n284_), .A4(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT93), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n282_), .A2(new_n284_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n293_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n294_), .A2(KEYINPUT21), .A3(new_n295_), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G228gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(new_n263_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  INV_X1    g102(.A(G141gat), .ZN(new_n304_));
  INV_X1    g103(.A(G148gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT1), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n303_), .B(new_n306_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G155gat), .B(G162gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT3), .ZN(new_n314_));
  AND3_X1   g113(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n313_), .A2(new_n314_), .B1(new_n315_), .B2(KEYINPUT86), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT87), .B(new_n311_), .C1(new_n316_), .C2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n314_), .A2(new_n313_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n318_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n317_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n311_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n322_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n310_), .B1(new_n321_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT88), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n332_), .B(new_n310_), .C1(new_n321_), .C2(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n302_), .B1(new_n334_), .B2(KEYINPUT29), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT94), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n292_), .A2(new_n297_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n301_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n280_), .B1(new_n335_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n327_), .A2(new_n328_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT87), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n327_), .A2(new_n322_), .A3(new_n328_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n344_), .B1(new_n348_), .B2(new_n310_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n298_), .A2(KEYINPUT94), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n337_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n300_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n344_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n352_), .B(new_n279_), .C1(new_n353_), .C2(new_n302_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n343_), .A2(KEYINPUT90), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G22gat), .B(G50gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n331_), .A2(new_n344_), .A3(new_n333_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n356_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n343_), .A2(new_n354_), .A3(KEYINPUT90), .A4(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n357_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n276_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n362_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n272_), .A2(new_n275_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n260_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n348_), .A2(new_n255_), .A3(new_n310_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT4), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n260_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n332_), .B1(new_n348_), .B2(new_n310_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n333_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT0), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G57gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n373_), .A2(new_n385_), .A3(new_n375_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n386_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n384_), .B1(new_n376_), .B2(new_n382_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n390_), .B1(new_n395_), .B2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT104), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT96), .B1(new_n238_), .B2(new_n224_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT25), .B(G183gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT26), .B(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n404_));
  INV_X1    g203(.A(new_n237_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n214_), .A2(new_n235_), .A3(KEYINPUT23), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n404_), .B(new_n225_), .C1(new_n407_), .C2(new_n234_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n400_), .A2(new_n223_), .A3(new_n403_), .A4(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n229_), .B1(new_n217_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n399_), .B1(new_n412_), .B2(new_n298_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n243_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n226_), .A2(new_n227_), .A3(new_n241_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n298_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT19), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n413_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT97), .B1(new_n412_), .B2(new_n298_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n298_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n409_), .A2(new_n416_), .A3(new_n424_), .A4(new_n411_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n423_), .A4(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n420_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT18), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G64gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G92gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n398_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n423_), .B(KEYINPUT20), .C1(new_n340_), .C2(new_n412_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n419_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n413_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT103), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT103), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n413_), .A2(new_n417_), .A3(new_n437_), .A4(new_n421_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n431_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n426_), .A2(new_n421_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n413_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n431_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT104), .A3(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n432_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT27), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n444_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n441_), .A2(new_n431_), .A3(new_n442_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT27), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n397_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n372_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n383_), .A2(new_n384_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n380_), .A2(new_n385_), .A3(new_n374_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n390_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT100), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n454_), .A2(KEYINPUT100), .A3(new_n390_), .A4(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n450_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n395_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(KEYINPUT33), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n394_), .A2(KEYINPUT99), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n386_), .A2(KEYINPUT33), .A3(new_n391_), .A4(new_n393_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT98), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n469_), .A3(KEYINPUT33), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n460_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n443_), .B1(new_n475_), .B2(new_n431_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n476_), .A2(KEYINPUT102), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n439_), .A2(KEYINPUT32), .A3(new_n444_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(KEYINPUT102), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n477_), .A2(new_n397_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n460_), .A2(new_n466_), .A3(new_n471_), .A4(KEYINPUT101), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n363_), .A2(new_n364_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(new_n276_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n453_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  INV_X1    g285(.A(G43gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G50gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G1gat), .ZN(new_n491_));
  INV_X1    g290(.A(G8gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT71), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G8gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n490_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n490_), .A2(new_n500_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n489_), .B(KEYINPUT15), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n500_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n504_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(new_n219_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(new_n281_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n508_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT78), .Z(new_n513_));
  INV_X1    g312(.A(KEYINPUT65), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n514_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  INV_X1    g315(.A(G99gat), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n278_), .A4(KEYINPUT65), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT6), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n515_), .B(new_n518_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  XOR2_X1   g323(.A(G85gat), .B(G92gat), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n525_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT67), .B1(new_n530_), .B2(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT67), .ZN(new_n532_));
  AOI211_X1 g331(.A(new_n532_), .B(new_n524_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n533_));
  OAI22_X1  g332(.A1(new_n528_), .A2(new_n529_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n525_), .A2(KEYINPUT9), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT10), .B(G99gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT64), .B(G106gat), .ZN(new_n539_));
  OAI221_X1 g338(.A(new_n536_), .B1(KEYINPUT9), .B2(new_n537_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n520_), .A2(new_n522_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n490_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT34), .Z(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n534_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n530_), .A2(KEYINPUT8), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n532_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n530_), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n526_), .B(new_n527_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(KEYINPUT68), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n542_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n544_), .B(new_n548_), .C1(new_n506_), .C2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n546_), .A2(new_n547_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G134gat), .ZN(new_n562_));
  INV_X1    g361(.A(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n560_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT69), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n560_), .A2(new_n566_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n560_), .A2(new_n571_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n569_), .A2(new_n570_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n568_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT37), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n500_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  NOR2_X1   g383(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n580_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(KEYINPUT17), .A3(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT75), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT76), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(new_n587_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n578_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n586_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n535_), .A2(new_n542_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n550_), .A2(new_n556_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n542_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n602_), .B1(new_n606_), .B2(new_n601_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n603_), .B1(new_n543_), .B2(new_n586_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n608_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n543_), .A2(new_n586_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n612_), .B2(new_n602_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G176gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n283_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(new_n613_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT13), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n600_), .A2(new_n623_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n485_), .B(new_n513_), .C1(new_n624_), .C2(KEYINPUT77), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(KEYINPUT77), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n397_), .B(KEYINPUT105), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n491_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT38), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n482_), .A2(new_n484_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n453_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n622_), .B(KEYINPUT13), .Z(new_n634_));
  INV_X1    g433(.A(new_n512_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n569_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n599_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n633_), .A2(new_n636_), .A3(new_n637_), .A4(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n397_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n630_), .A2(new_n641_), .ZN(G1324gat));
  NAND2_X1  g441(.A1(new_n447_), .A2(new_n451_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G8gat), .B1(new_n639_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT106), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n646_), .B(G8gat), .C1(new_n639_), .C2(new_n643_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(KEYINPUT39), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n643_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n625_), .A2(new_n492_), .A3(new_n649_), .A4(new_n626_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(KEYINPUT106), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT107), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n648_), .A2(new_n655_), .A3(new_n650_), .A4(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  OAI21_X1  g458(.A(G15gat), .B1(new_n639_), .B2(new_n369_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT41), .Z(new_n661_));
  INV_X1    g460(.A(G15gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n627_), .A2(new_n662_), .A3(new_n276_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n627_), .A2(new_n665_), .A3(new_n483_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n483_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n639_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT108), .Z(G1327gat));
  INV_X1    g470(.A(new_n513_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n638_), .A2(new_n637_), .ZN(new_n673_));
  AND4_X1   g472(.A1(new_n623_), .A2(new_n633_), .A3(new_n672_), .A4(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(G29gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n397_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n628_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n633_), .A2(KEYINPUT43), .A3(new_n578_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(new_n485_), .B2(new_n577_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(KEYINPUT109), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n635_), .B(new_n634_), .C1(KEYINPUT109), .C2(new_n682_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n681_), .A2(new_n599_), .A3(new_n684_), .A4(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n678_), .A2(new_n680_), .A3(new_n599_), .A4(new_n685_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n683_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n677_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n676_), .B1(new_n689_), .B2(new_n675_), .ZN(G1328gat));
  AND2_X1   g489(.A1(new_n687_), .A2(new_n683_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n687_), .A2(new_n683_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n649_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT110), .B(new_n649_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(G36gat), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT111), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT112), .Z(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n674_), .A2(new_n701_), .A3(new_n649_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT45), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n697_), .A2(new_n700_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n700_), .B1(new_n697_), .B2(new_n703_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND2_X1  g505(.A1(new_n674_), .A2(new_n276_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT114), .B(G43gat), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n487_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n710_), .A2(KEYINPUT113), .A3(new_n276_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT113), .B1(new_n710_), .B2(new_n276_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n709_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  INV_X1    g516(.A(G50gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n674_), .A2(new_n718_), .A3(new_n483_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n667_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n718_), .ZN(G1331gat));
  NOR3_X1   g520(.A1(new_n485_), .A2(new_n512_), .A3(new_n623_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n600_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT115), .Z(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n628_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n637_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n485_), .A2(new_n726_), .A3(new_n599_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n634_), .A3(new_n513_), .ZN(new_n728_));
  INV_X1    g527(.A(G57gat), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n640_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT116), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n725_), .A2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n733_), .A3(new_n649_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G64gat), .B1(new_n728_), .B2(new_n643_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT48), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n738_), .A3(new_n276_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G71gat), .B1(new_n728_), .B2(new_n369_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT49), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n724_), .A2(new_n743_), .A3(new_n483_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G78gat), .B1(new_n728_), .B2(new_n667_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1335gat));
  AND2_X1   g546(.A1(new_n722_), .A2(new_n673_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n628_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n623_), .A2(new_n512_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n678_), .A2(new_n680_), .A3(new_n599_), .A4(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n397_), .A2(G85gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  AOI21_X1  g553(.A(G92gat), .B1(new_n748_), .B2(new_n649_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n649_), .A2(G92gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n752_), .B2(new_n756_), .ZN(G1337gat));
  OAI21_X1  g556(.A(G99gat), .B1(new_n751_), .B2(new_n369_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n538_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n748_), .A2(new_n761_), .A3(new_n276_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n759_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(KEYINPUT118), .B2(KEYINPUT51), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n765_), .A2(new_n768_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n764_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1338gat));
  OAI21_X1  g570(.A(G106gat), .B1(new_n751_), .B2(new_n667_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT52), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(G106gat), .C1(new_n751_), .C2(new_n667_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n667_), .A2(new_n539_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n748_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT119), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n776_), .A2(new_n781_), .A3(new_n778_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT53), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n778_), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT119), .B(new_n785_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n784_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n783_), .A2(new_n788_), .ZN(G1339gat));
  NOR2_X1   g588(.A1(new_n649_), .A2(new_n365_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n608_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n610_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n534_), .A2(new_n549_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT68), .B1(new_n554_), .B2(new_n555_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n605_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT12), .A3(new_n601_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n602_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n609_), .A3(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n800_), .A2(new_n793_), .A3(new_n611_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n620_), .B1(new_n794_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n791_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n512_), .A2(new_n621_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n793_), .B1(new_n800_), .B2(new_n611_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n800_), .A2(new_n611_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n618_), .B1(new_n809_), .B2(new_n801_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n806_), .A3(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n508_), .A2(new_n511_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n501_), .A2(new_n502_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(new_n511_), .C1(new_n502_), .C2(new_n507_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n622_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT57), .B1(new_n817_), .B2(new_n637_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n819_), .B(new_n726_), .C1(new_n812_), .C2(new_n816_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n813_), .A2(new_n815_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n810_), .B2(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n803_), .A2(new_n791_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n621_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n621_), .A4(new_n824_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n578_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n638_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n577_), .A2(new_n623_), .A3(new_n638_), .A4(new_n513_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT54), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n628_), .B(new_n790_), .C1(new_n830_), .C2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n512_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n827_), .A2(new_n578_), .A3(new_n828_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n839_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n832_), .B1(new_n840_), .B2(new_n638_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n628_), .A4(new_n790_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n838_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(G113gat), .A3(new_n672_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n835_), .A2(new_n512_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(KEYINPUT121), .A3(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n837_), .A2(new_n845_), .A3(new_n848_), .ZN(G1340gat));
  NAND3_X1  g648(.A1(new_n838_), .A2(new_n634_), .A3(new_n843_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G120gat), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n623_), .B2(G120gat), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n835_), .B(new_n853_), .C1(new_n852_), .C2(G120gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT122), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n851_), .A2(new_n854_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n835_), .B2(new_n638_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n638_), .A2(G127gat), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT123), .Z(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n844_), .B2(new_n862_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n835_), .B2(new_n726_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n578_), .A2(G134gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n844_), .B2(new_n865_), .ZN(G1343gat));
  INV_X1    g665(.A(new_n371_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n841_), .A2(new_n867_), .A3(new_n643_), .A4(new_n628_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n635_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n304_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n623_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n305_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n599_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT124), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n873_), .B(new_n875_), .ZN(G1346gat));
  NOR3_X1   g675(.A1(new_n868_), .A2(new_n563_), .A3(new_n577_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n563_), .B1(new_n868_), .B2(new_n637_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n879_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n880_), .B2(new_n881_), .ZN(G1347gat));
  NAND2_X1  g681(.A1(new_n821_), .A2(new_n829_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n599_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n643_), .B1(new_n884_), .B2(new_n832_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n628_), .A2(new_n365_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n885_), .A2(KEYINPUT126), .A3(new_n512_), .A4(new_n886_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n841_), .A2(new_n512_), .A3(new_n649_), .A4(new_n886_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(G169gat), .A3(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n891_), .A2(KEYINPUT62), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n885_), .A2(new_n886_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT22), .B(G169gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n512_), .A2(new_n895_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT127), .Z(new_n897_));
  OAI22_X1  g696(.A1(new_n892_), .A2(new_n893_), .B1(new_n894_), .B2(new_n897_), .ZN(G1348gat));
  NOR2_X1   g697(.A1(new_n894_), .A2(new_n623_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n220_), .ZN(G1349gat));
  INV_X1    g699(.A(new_n894_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n638_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n401_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n239_), .B2(new_n902_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n894_), .B2(new_n577_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n726_), .A2(new_n402_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n894_), .B2(new_n906_), .ZN(G1351gat));
  AND3_X1   g706(.A1(new_n841_), .A2(new_n640_), .A3(new_n649_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n867_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n635_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n281_), .ZN(G1352gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n623_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n283_), .ZN(G1353gat));
  INV_X1    g712(.A(new_n909_), .ZN(new_n914_));
  AOI211_X1 g713(.A(KEYINPUT63), .B(G211gat), .C1(new_n914_), .C2(new_n638_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT63), .B(G211gat), .Z(new_n916_));
  AND3_X1   g715(.A1(new_n914_), .A2(new_n638_), .A3(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1354gat));
  AND3_X1   g717(.A1(new_n914_), .A2(G218gat), .A3(new_n578_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n914_), .B2(new_n726_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1355gat));
endmodule


