//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT66), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(KEYINPUT65), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n209_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n202_), .B1(new_n208_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n218_), .B(new_n202_), .C1(new_n213_), .C2(new_n207_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n214_), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G57gat), .B(G64gat), .Z(new_n222_));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT68), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n222_), .A2(new_n223_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n227_), .A2(KEYINPUT68), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(KEYINPUT68), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT10), .B(G99gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT9), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G85gat), .A3(G92gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n207_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n221_), .A2(new_n235_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n235_), .B1(new_n221_), .B2(new_n243_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(KEYINPUT69), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n221_), .A2(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n235_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT70), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n221_), .A2(new_n243_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n235_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT12), .A3(new_n244_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n251_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n250_), .A2(new_n263_), .A3(new_n252_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G120gat), .B(G148gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n254_), .A2(new_n262_), .A3(new_n264_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT72), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n263_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n273_));
  AOI211_X1 g072(.A(KEYINPUT70), .B(new_n251_), .C1(new_n246_), .C2(new_n249_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n262_), .A4(new_n270_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n262_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n269_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT13), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n286_));
  INV_X1    g085(.A(G197gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G204gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT88), .B1(new_n285_), .B2(G197gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT21), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(G197gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n288_), .A4(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n288_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT21), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n300_), .B2(new_n296_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n296_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n302_), .A2(KEYINPUT90), .A3(KEYINPUT21), .A4(new_n299_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306_));
  INV_X1    g105(.A(G190gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(KEYINPUT26), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n305_), .B(new_n308_), .C1(new_n309_), .C2(new_n306_), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n310_), .A2(KEYINPUT79), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT79), .B1(new_n310_), .B2(new_n315_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n319_), .A2(new_n322_), .A3(KEYINPUT80), .A4(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n316_), .A2(new_n317_), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT81), .B1(new_n311_), .B2(KEYINPUT22), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n312_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332_));
  XOR2_X1   g131(.A(KEYINPUT22), .B(G169gat), .Z(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n322_), .B(new_n323_), .C1(G183gat), .C2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n314_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n304_), .B1(new_n329_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n309_), .A2(new_n305_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n315_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n333_), .A2(G176gat), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n340_), .A2(new_n324_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n304_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(KEYINPUT20), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT94), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G64gat), .ZN(new_n352_));
  INV_X1    g151(.A(G92gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n304_), .A2(new_n342_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT95), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT95), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n304_), .A2(new_n358_), .A3(new_n342_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n310_), .A2(new_n315_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n310_), .A2(KEYINPUT79), .A3(new_n315_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n328_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n304_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n337_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n360_), .A2(KEYINPUT20), .A3(new_n347_), .A4(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n349_), .A2(new_n355_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n355_), .B1(new_n349_), .B2(new_n370_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n284_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n359_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n358_), .B1(new_n304_), .B2(new_n342_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n369_), .B(KEYINPUT20), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n348_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n366_), .A2(new_n368_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n304_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n347_), .B1(new_n382_), .B2(new_n343_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n354_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n349_), .A2(new_n355_), .A3(new_n370_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT98), .A3(new_n284_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n375_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n378_), .A2(new_n347_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n348_), .B1(new_n382_), .B2(new_n343_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n355_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(new_n391_), .A3(KEYINPUT27), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  INV_X1    g195(.A(G155gat), .ZN(new_n397_));
  INV_X1    g196(.A(G162gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT1), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT1), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G155gat), .A3(G162gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n399_), .B(new_n401_), .C1(G155gat), .C2(G162gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G141gat), .ZN(new_n408_));
  INV_X1    g207(.A(G148gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n402_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT2), .B1(new_n405_), .B2(new_n406_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT2), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n403_), .A2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n412_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n397_), .A2(new_n398_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n411_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G127gat), .A2(G134gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G127gat), .A2(G134gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n425_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G127gat), .ZN(new_n430_));
  INV_X1    g229(.A(G134gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT84), .A3(new_n426_), .ZN(new_n433_));
  AND2_X1   g232(.A1(G113gat), .A2(G120gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G113gat), .A2(G120gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n429_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT85), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(KEYINPUT85), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n424_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n406_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n417_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n418_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n415_), .A4(new_n414_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n407_), .A2(new_n410_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n446_), .A2(new_n422_), .B1(new_n447_), .B2(new_n402_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n429_), .A2(new_n433_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n436_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n429_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n396_), .B1(new_n441_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n438_), .A2(KEYINPUT85), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n453_), .B2(KEYINPUT85), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT4), .B1(new_n457_), .B2(new_n424_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n395_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(G85gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT0), .ZN(new_n462_));
  INV_X1    g261(.A(G57gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n441_), .A2(new_n394_), .A3(new_n454_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n464_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G50gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT28), .B1(new_n424_), .B2(KEYINPUT29), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT28), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n448_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G22gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n470_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G22gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G50gat), .A3(new_n476_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT87), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n448_), .A2(new_n473_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(new_n367_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G78gat), .B(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n424_), .A2(KEYINPUT29), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n304_), .A3(new_n485_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n488_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n489_), .B(KEYINPUT91), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n485_), .B1(new_n490_), .B2(new_n304_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n483_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n488_), .A2(new_n491_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n494_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n488_), .A2(new_n493_), .A3(new_n491_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n502_), .A2(new_n503_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n503_), .A2(KEYINPUT92), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n497_), .A2(KEYINPUT92), .A3(new_n503_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n483_), .A2(new_n508_), .A3(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT93), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n499_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT82), .B(KEYINPUT30), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n457_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(new_n381_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT83), .B(G99gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT31), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G43gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G71gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n514_), .B(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n393_), .A2(new_n469_), .A3(new_n511_), .A4(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n499_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n505_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n526_));
  AND4_X1   g325(.A1(new_n505_), .A2(new_n483_), .A3(new_n508_), .A4(new_n506_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n388_), .A2(new_n469_), .A3(new_n528_), .A4(new_n392_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n466_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n466_), .B2(new_n530_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n441_), .A2(new_n454_), .A3(new_n395_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n455_), .A2(new_n458_), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n464_), .B(new_n534_), .C1(new_n535_), .C2(new_n394_), .ZN(new_n536_));
  NOR4_X1   g335(.A1(new_n386_), .A2(new_n532_), .A3(new_n533_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n538_), .B(new_n539_), .C1(new_n379_), .C2(new_n383_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT32), .B(new_n354_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n349_), .A2(new_n370_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n543_), .B2(new_n539_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n542_), .A2(new_n544_), .A3(new_n469_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n511_), .B1(new_n537_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n529_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n522_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT99), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT99), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n551_), .A3(new_n548_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n524_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G29gat), .B(G36gat), .ZN(new_n554_));
  INV_X1    g353(.A(G43gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n470_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT15), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559_));
  INV_X1    g358(.A(G1gat), .ZN(new_n560_));
  INV_X1    g359(.A(G8gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G1gat), .B(G8gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n557_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n558_), .A2(KEYINPUT75), .A3(new_n565_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n568_), .A2(new_n569_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n557_), .B(new_n570_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n311_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n287_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n573_), .A2(new_n576_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(KEYINPUT76), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n585_), .A3(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT77), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n283_), .A2(new_n553_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n255_), .A2(new_n558_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT73), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n247_), .A2(new_n557_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n594_), .A2(new_n595_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n591_), .A2(KEYINPUT35), .A3(new_n593_), .A4(new_n597_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G134gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n398_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n601_), .A2(new_n602_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n606_), .B(KEYINPUT36), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n601_), .A2(new_n611_), .A3(new_n602_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n608_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT37), .B1(new_n614_), .B2(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n565_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n235_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(G183gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(G211gat), .Z(new_n624_));
  NOR3_X1   g423(.A1(new_n619_), .A2(new_n620_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(KEYINPUT17), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n616_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT74), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n589_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n469_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n560_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT38), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n608_), .A2(new_n612_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT100), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n553_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n283_), .A2(new_n587_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n627_), .A3(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT101), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT101), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n633_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT102), .A3(G1gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT102), .B1(new_n645_), .B2(G1gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n635_), .B1(new_n646_), .B2(new_n647_), .ZN(G1324gat));
  OAI21_X1  g447(.A(G8gat), .B1(new_n641_), .B2(new_n393_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(G8gat), .C1(new_n641_), .C2(new_n393_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n393_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n632_), .A2(new_n561_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT103), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n653_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n657_), .A2(KEYINPUT40), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT40), .B1(new_n657_), .B2(new_n659_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OR3_X1    g461(.A1(new_n631_), .A2(G15gat), .A3(new_n548_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n642_), .A2(new_n522_), .A3(new_n643_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT41), .B1(new_n664_), .B2(G15gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT104), .B(new_n663_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1326gat));
  NAND3_X1  g470(.A1(new_n632_), .A2(new_n475_), .A3(new_n528_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n644_), .A2(new_n528_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(G22gat), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT42), .B(new_n475_), .C1(new_n644_), .C2(new_n528_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(new_n587_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n281_), .A2(KEYINPUT13), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT13), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n628_), .B(new_n678_), .C1(new_n679_), .C2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n616_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n553_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n551_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT99), .B(new_n522_), .C1(new_n529_), .C2(new_n546_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n523_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n616_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n682_), .B1(new_n684_), .B2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT106), .B1(new_n690_), .B2(KEYINPUT105), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  INV_X1    g491(.A(new_n682_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n687_), .A2(new_n688_), .A3(new_n616_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n688_), .B1(new_n687_), .B2(new_n616_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n692_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n691_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT106), .B(new_n692_), .C1(new_n690_), .C2(KEYINPUT105), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n469_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n588_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n636_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n627_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n282_), .A2(new_n687_), .A3(new_n704_), .A4(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT107), .Z(new_n708_));
  INV_X1    g507(.A(G29gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n633_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n703_), .A2(new_n710_), .ZN(G1328gat));
  XNOR2_X1  g510(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT108), .B1(new_n701_), .B2(new_n654_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n715_), .B(new_n393_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n714_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n708_), .A2(new_n717_), .A3(new_n654_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n713_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n714_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n716_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n720_), .A3(new_n712_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n726_), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n708_), .A2(new_n555_), .A3(new_n522_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n548_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n555_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT110), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n728_), .B(new_n732_), .C1(new_n729_), .C2(new_n555_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n731_), .A2(KEYINPUT47), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT47), .B1(new_n731_), .B2(new_n733_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1330gat));
  OAI21_X1  g535(.A(G50gat), .B1(new_n702_), .B2(new_n511_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n708_), .A2(new_n470_), .A3(new_n528_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n282_), .A2(new_n553_), .A3(new_n678_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n630_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n633_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT111), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n639_), .A2(new_n627_), .A3(new_n283_), .A4(new_n588_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n633_), .A2(G57gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT112), .ZN(G1332gat));
  OAI21_X1  g546(.A(G64gat), .B1(new_n744_), .B2(new_n393_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  INV_X1    g548(.A(new_n741_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n393_), .A2(G64gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT113), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n744_), .B2(new_n548_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n548_), .A2(G71gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n750_), .B2(new_n756_), .ZN(G1334gat));
  OAI21_X1  g556(.A(G78gat), .B1(new_n744_), .B2(new_n511_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT50), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n511_), .A2(G78gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n750_), .B2(new_n760_), .ZN(G1335gat));
  AND2_X1   g560(.A1(new_n740_), .A2(new_n706_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n633_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n684_), .A2(new_n689_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n282_), .A2(new_n678_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n628_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n633_), .A2(G85gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n766_), .B2(new_n393_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n762_), .A2(new_n353_), .A3(new_n654_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT114), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n522_), .A3(new_n236_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n764_), .A2(new_n628_), .A3(new_n522_), .A4(new_n765_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT115), .B1(new_n775_), .B2(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT116), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(KEYINPUT116), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(KEYINPUT51), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT51), .B1(new_n780_), .B2(new_n781_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n766_), .B2(new_n511_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT118), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(G106gat), .C1(new_n766_), .C2(new_n511_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n762_), .A2(new_n528_), .A3(new_n237_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT117), .Z(new_n793_));
  NAND3_X1  g592(.A1(new_n786_), .A2(KEYINPUT52), .A3(new_n788_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n282_), .A2(new_n629_), .A3(new_n588_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT119), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n282_), .A2(new_n629_), .A3(new_n799_), .A4(new_n588_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n798_), .A2(KEYINPUT54), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT54), .B1(new_n798_), .B2(new_n800_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n568_), .A2(new_n575_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n574_), .A2(new_n569_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n580_), .A3(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n583_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n281_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT120), .B1(new_n278_), .B2(new_n678_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n811_), .B(new_n587_), .C1(new_n272_), .C2(new_n277_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n258_), .A2(new_n252_), .A3(new_n260_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT121), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n258_), .A2(new_n816_), .A3(new_n252_), .A4(new_n260_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(new_n261_), .B2(new_n251_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n252_), .C1(new_n258_), .C2(new_n260_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n270_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT122), .B1(new_n823_), .B2(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n262_), .A2(new_n820_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n261_), .A2(KEYINPUT55), .A3(new_n251_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n815_), .A3(new_n817_), .A4(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n269_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n828_), .A2(new_n830_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n809_), .B1(new_n813_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n804_), .B1(new_n836_), .B2(new_n636_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n833_), .B1(new_n824_), .B2(new_n831_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n838_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT57), .B(new_n705_), .C1(new_n839_), .C2(new_n809_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n823_), .A2(KEYINPUT56), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n278_), .B(new_n808_), .C1(new_n833_), .C2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n843_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n616_), .A3(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n837_), .A2(new_n840_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n628_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n803_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n654_), .A2(new_n469_), .A3(new_n528_), .A4(new_n548_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n704_), .A2(G113gat), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n847_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n837_), .A2(new_n840_), .A3(new_n846_), .A4(KEYINPUT123), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n628_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n803_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n858_), .A2(new_n851_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n852_), .B(new_n853_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G113gat), .B1(new_n859_), .B2(new_n678_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1340gat));
  OAI211_X1 g662(.A(new_n283_), .B(new_n852_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT124), .B(G120gat), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n282_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n859_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n867_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n869_), .ZN(G1341gat));
  NOR2_X1   g669(.A1(new_n628_), .A2(new_n430_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n852_), .B(new_n871_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G127gat), .B1(new_n859_), .B2(new_n627_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  NOR2_X1   g674(.A1(new_n683_), .A2(new_n431_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n852_), .B(new_n876_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G134gat), .B1(new_n859_), .B2(new_n638_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n511_), .A2(new_n522_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n857_), .B2(new_n803_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n883_), .A2(new_n633_), .A3(new_n393_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n678_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G141gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n408_), .A3(new_n678_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n283_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G148gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n884_), .A2(new_n409_), .A3(new_n283_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1345gat));
  NAND2_X1  g691(.A1(new_n884_), .A2(new_n627_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT125), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n884_), .A2(new_n627_), .A3(new_n895_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1346gat));
  NAND2_X1  g698(.A1(new_n884_), .A2(new_n638_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n683_), .A2(new_n398_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n900_), .A2(new_n398_), .B1(new_n884_), .B2(new_n901_), .ZN(G1347gat));
  NOR4_X1   g701(.A1(new_n393_), .A2(new_n633_), .A3(new_n528_), .A4(new_n548_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n849_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n678_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n587_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n311_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n907_), .B(new_n910_), .C1(new_n333_), .C2(new_n906_), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n905_), .B2(new_n283_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n312_), .B(new_n282_), .C1(new_n857_), .C2(new_n803_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n913_), .ZN(G1349gat));
  NOR2_X1   g713(.A1(new_n904_), .A2(new_n628_), .ZN(new_n915_));
  MUX2_X1   g714(.A(G183gat), .B(new_n305_), .S(new_n915_), .Z(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n904_), .B2(new_n683_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n638_), .A2(new_n309_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n904_), .B2(new_n918_), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n393_), .A2(new_n633_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n883_), .A2(new_n678_), .A3(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g721(.A1(new_n883_), .A2(new_n920_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n283_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G204gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n285_), .A3(new_n283_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n883_), .A2(new_n627_), .A3(new_n920_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AND2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n928_), .B2(new_n929_), .ZN(G1354gat));
  NAND4_X1  g731(.A1(new_n858_), .A2(new_n638_), .A3(new_n881_), .A4(new_n920_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(G218gat), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n883_), .A2(KEYINPUT126), .A3(new_n638_), .A4(new_n920_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n616_), .A2(G218gat), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(KEYINPUT127), .Z(new_n940_));
  NAND2_X1  g739(.A1(new_n923_), .A2(new_n940_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n938_), .A2(new_n941_), .ZN(G1355gat));
endmodule


