//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n202_));
  INV_X1    g001(.A(G71gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT66), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G71gat), .ZN(new_n206_));
  INV_X1    g005(.A(G78gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n202_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(G71gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n203_), .A2(KEYINPUT66), .ZN(new_n212_));
  OAI21_X1  g011(.A(G78gat), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT11), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G57gat), .B(G64gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n216_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT11), .A4(new_n214_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n223_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G85gat), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT64), .A3(new_n224_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  INV_X1    g038(.A(G99gat), .ZN(new_n240_));
  INV_X1    g039(.A(G106gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n236_), .A2(new_n237_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n243_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(KEYINPUT65), .A3(new_n243_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n232_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n246_), .B1(new_n252_), .B2(new_n245_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n254_));
  OR2_X1    g053(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n241_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n230_), .A2(KEYINPUT9), .A3(new_n224_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n238_), .A2(new_n254_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n217_), .A2(KEYINPUT67), .A3(new_n219_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n222_), .A2(new_n253_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n217_), .A2(KEYINPUT67), .A3(new_n219_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT67), .B1(new_n217_), .B2(new_n219_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n243_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n249_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n251_), .A3(new_n238_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n245_), .B1(new_n270_), .B2(new_n233_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n248_), .A2(new_n247_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n272_), .A2(new_n232_), .A3(KEYINPUT8), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n259_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n275_), .A3(KEYINPUT68), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n263_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G230gat), .ZN(new_n279_));
  INV_X1    g078(.A(G233gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n217_), .A2(KEYINPUT12), .A3(new_n219_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n259_), .B(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n253_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n277_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n281_), .B1(new_n266_), .B2(new_n275_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G120gat), .B(G148gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G176gat), .B(G204gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n291_), .A2(new_n297_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT13), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT13), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n298_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n305_), .A2(KEYINPUT71), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(KEYINPUT71), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G8gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT76), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(KEYINPUT76), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G15gat), .B(G22gat), .ZN(new_n314_));
  INV_X1    g113(.A(G1gat), .ZN(new_n315_));
  INV_X1    g114(.A(G8gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT14), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n311_), .A2(new_n317_), .A3(new_n314_), .A4(new_n312_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G43gat), .B(G50gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G36gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G29gat), .ZN(new_n325_));
  INV_X1    g124(.A(G29gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G36gat), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT73), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT73), .B1(new_n325_), .B2(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n323_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n326_), .A2(G36gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n324_), .A2(G29gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT73), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n322_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n321_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n321_), .A2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n309_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT80), .A3(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G229gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT15), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n337_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n330_), .A2(new_n336_), .A3(KEYINPUT15), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(new_n321_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n344_), .A3(new_n338_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G113gat), .B(G141gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(G169gat), .B(G197gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n308_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT1), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n364_), .B(new_n366_), .C1(KEYINPUT1), .C2(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n370_), .B(KEYINPUT3), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n368_), .B(KEYINPUT2), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n366_), .A2(new_n361_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT85), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G120gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n382_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n367_), .A2(new_n371_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n386_), .A2(new_n388_), .A3(KEYINPUT4), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n378_), .A2(new_n394_), .A3(new_n385_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n390_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G1gat), .B(G29gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT95), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  OR3_X1    g200(.A1(new_n392_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  INV_X1    g209(.A(G169gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n411_), .A2(KEYINPUT22), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n412_), .B2(KEYINPUT81), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n406_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT23), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(G183gat), .B2(G190gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n415_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n411_), .A2(new_n410_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT24), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT24), .A3(new_n406_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n418_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT26), .B(G190gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT25), .B(G183gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n421_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G197gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G204gat), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n432_), .A2(KEYINPUT88), .ZN(new_n433_));
  INV_X1    g232(.A(G204gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G197gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(KEYINPUT88), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G211gat), .B(G218gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT21), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n435_), .B2(new_n432_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT87), .Z(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n437_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n441_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n430_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G226gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT19), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n427_), .B(KEYINPUT92), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n426_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n425_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n407_), .A2(new_n410_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n419_), .A2(new_n406_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT20), .B1(new_n455_), .B2(new_n446_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n447_), .A2(new_n449_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n430_), .A2(new_n446_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n446_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT93), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n457_), .B1(new_n463_), .B2(new_n449_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G8gat), .B(G36gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n449_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n473_), .B2(new_n457_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT27), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n456_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n447_), .B1(KEYINPUT98), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(KEYINPUT98), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n472_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n463_), .A2(new_n449_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n471_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n475_), .A2(new_n476_), .B1(new_n477_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n385_), .B(KEYINPUT31), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n430_), .B(KEYINPUT30), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT83), .B(G43gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n430_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G71gat), .B(G99gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT84), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G15gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n491_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n488_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n493_), .A2(new_n494_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n489_), .A2(new_n490_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n498_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n487_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT91), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n378_), .A2(KEYINPUT29), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n446_), .ZN(new_n512_));
  INV_X1    g311(.A(G228gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(new_n280_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n512_), .A2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n510_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G22gat), .B(G50gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT29), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n387_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n520_), .B1(new_n387_), .B2(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n522_), .A3(new_n518_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n512_), .A2(new_n514_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n511_), .B(new_n446_), .C1(new_n513_), .C2(new_n280_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n530_), .B(new_n531_), .C1(KEYINPUT91), .C2(new_n509_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n517_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n508_), .B(KEYINPUT90), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n509_), .A2(KEYINPUT90), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n537_), .A3(new_n528_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n533_), .A2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n502_), .A2(new_n507_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n405_), .B(new_n484_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n469_), .A2(KEYINPUT32), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n464_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n481_), .A2(new_n482_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n404_), .B(new_n544_), .C1(new_n545_), .C2(new_n543_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n403_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT97), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n401_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n393_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(KEYINPUT33), .B(new_n401_), .C1(new_n392_), .C2(new_n396_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n470_), .A2(new_n474_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n546_), .B1(new_n549_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n539_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n542_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n360_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT74), .ZN(new_n562_));
  XOR2_X1   g361(.A(G134gat), .B(G162gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n350_), .B1(new_n253_), .B2(new_n285_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n337_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n274_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n350_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n253_), .A2(new_n285_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n571_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n253_), .A2(new_n337_), .A3(new_n259_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n573_), .A4(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n566_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n565_), .B1(new_n583_), .B2(new_n564_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n576_), .A2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT75), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n586_), .B(new_n565_), .C1(new_n583_), .C2(new_n564_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n588_), .A2(KEYINPUT37), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT37), .B1(new_n588_), .B2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT17), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT78), .ZN(new_n598_));
  AND2_X1   g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n321_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n266_), .A2(KEYINPUT77), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n266_), .A2(KEYINPUT77), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n600_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n601_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n220_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n600_), .A2(new_n220_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n596_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n592_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT79), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n560_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n404_), .A2(new_n315_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n308_), .A2(new_n615_), .A3(new_n359_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n588_), .A2(new_n589_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n559_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT100), .B1(new_n559_), .B2(new_n625_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n405_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n623_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT101), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n623_), .A2(new_n634_), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(new_n619_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n484_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n316_), .A3(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n624_), .B(new_n638_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G8gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT102), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n640_), .A2(new_n644_), .A3(G8gat), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n642_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n643_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n639_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT40), .B(new_n639_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1325gat));
  NAND2_X1  g451(.A1(new_n502_), .A2(new_n507_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G15gat), .B1(new_n630_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n619_), .A2(G15gat), .A3(new_n653_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  OAI21_X1  g456(.A(G22gat), .B1(new_n630_), .B2(new_n539_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n658_), .B(new_n659_), .Z(new_n660_));
  NOR3_X1   g459(.A1(new_n619_), .A2(G22gat), .A3(new_n539_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n625_), .A2(new_n616_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n360_), .A2(new_n559_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n404_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n308_), .A2(new_n616_), .A3(new_n359_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  INV_X1    g467(.A(new_n591_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n588_), .A2(KEYINPUT37), .A3(new_n589_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n559_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n559_), .B2(new_n671_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT104), .B(new_n668_), .C1(new_n559_), .C2(new_n671_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n667_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n678_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n667_), .B(new_n681_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n405_), .A2(new_n326_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n666_), .B1(new_n684_), .B2(new_n685_), .ZN(G1328gat));
  XNOR2_X1  g485(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n484_), .A2(G36gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n664_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n664_), .B2(new_n689_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n679_), .A2(new_n682_), .A3(new_n638_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G36gat), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n694_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1329gat));
  INV_X1    g500(.A(new_n653_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n679_), .A2(new_n682_), .A3(G43gat), .A4(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n664_), .A2(new_n653_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(G43gat), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g505(.A1(new_n680_), .A2(new_n539_), .A3(new_n683_), .ZN(new_n707_));
  INV_X1    g506(.A(G50gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n556_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT108), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n707_), .A2(new_n708_), .B1(new_n664_), .B2(new_n710_), .ZN(G1331gat));
  NAND2_X1  g510(.A1(new_n618_), .A2(new_n308_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(KEYINPUT109), .ZN(new_n713_));
  INV_X1    g512(.A(new_n359_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n542_), .B2(new_n558_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(KEYINPUT109), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n404_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n308_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n616_), .A2(new_n359_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n628_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n629_), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n719_), .B(new_n720_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n404_), .B2(KEYINPUT110), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(KEYINPUT110), .B2(new_n724_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n718_), .B1(new_n723_), .B2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n723_), .B2(new_n638_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT48), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n717_), .A2(new_n728_), .A3(new_n638_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1333gat));
  AOI21_X1  g531(.A(new_n203_), .B1(new_n723_), .B2(new_n702_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n717_), .A2(new_n203_), .A3(new_n702_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1334gat));
  AOI21_X1  g535(.A(new_n207_), .B1(new_n723_), .B2(new_n556_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT50), .Z(new_n738_));
  NAND2_X1  g537(.A1(new_n556_), .A2(new_n207_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n717_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1335gat));
  AND3_X1   g541(.A1(new_n308_), .A2(new_n715_), .A3(new_n663_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n404_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n675_), .A2(new_n676_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n719_), .A2(new_n616_), .A3(new_n714_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(KEYINPUT112), .A3(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n405_), .A2(new_n228_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n744_), .B1(new_n753_), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n743_), .B2(new_n638_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n484_), .A2(new_n229_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n753_), .B2(new_n757_), .ZN(G1337gat));
  NAND4_X1  g557(.A1(new_n743_), .A2(new_n255_), .A3(new_n256_), .A4(new_n702_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n653_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n240_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(KEYINPUT51), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT51), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n759_), .C1(new_n760_), .C2(new_n240_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n743_), .A2(new_n241_), .A3(new_n556_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n745_), .A2(new_n556_), .A3(new_n746_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n339_), .A2(new_n344_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n355_), .B1(new_n779_), .B2(new_n351_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n356_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n302_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n286_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n222_), .A2(new_n260_), .B1(new_n253_), .B2(new_n259_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(KEYINPUT12), .ZN(new_n786_));
  INV_X1    g585(.A(new_n261_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n281_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n288_), .A2(new_n789_), .A3(new_n289_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n297_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n296_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT117), .B1(new_n792_), .B2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n792_), .A2(KEYINPUT117), .A3(new_n795_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n783_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n777_), .B(new_n671_), .C1(new_n799_), .C2(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(KEYINPUT58), .ZN(new_n801_));
  INV_X1    g600(.A(new_n281_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n288_), .B2(new_n261_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n261_), .A2(new_n802_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT55), .B1(new_n786_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n288_), .A2(new_n789_), .A3(new_n289_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n803_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n794_), .B1(new_n807_), .B2(new_n296_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  INV_X1    g608(.A(new_n795_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n807_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n811_), .A3(new_n798_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n782_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n300_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT58), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(new_n815_), .B2(new_n592_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n800_), .A2(new_n801_), .A3(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n807_), .A2(new_n810_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n714_), .B(new_n302_), .C1(new_n793_), .C2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n782_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n625_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  INV_X1    g622(.A(new_n625_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n823_), .B(new_n824_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n616_), .B1(new_n817_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n720_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(new_n592_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n828_), .B2(new_n592_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n827_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n540_), .A2(new_n484_), .A3(new_n404_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n833_), .A2(KEYINPUT59), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n822_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(KEYINPUT116), .B2(new_n825_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n821_), .A2(new_n625_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n823_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n817_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n832_), .B1(new_n843_), .B2(new_n615_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n834_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n835_), .A2(new_n836_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n837_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847_), .B2(new_n359_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n844_), .A2(new_n834_), .ZN(new_n849_));
  INV_X1    g648(.A(G113gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n714_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1340gat));
  OAI21_X1  g651(.A(G120gat), .B1(new_n847_), .B2(new_n719_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n719_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n849_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT120), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1341gat));
  OAI21_X1  g657(.A(G127gat), .B1(new_n847_), .B2(new_n615_), .ZN(new_n859_));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n849_), .A2(new_n860_), .A3(new_n616_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1342gat));
  OAI21_X1  g661(.A(G134gat), .B1(new_n847_), .B2(new_n592_), .ZN(new_n863_));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n849_), .A2(new_n864_), .A3(new_n824_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1343gat));
  INV_X1    g665(.A(new_n844_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n484_), .A2(new_n541_), .A3(new_n404_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n714_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n719_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(G148gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n616_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  OR3_X1    g677(.A1(new_n869_), .A2(G162gat), .A3(new_n625_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G162gat), .B1(new_n869_), .B2(new_n592_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n638_), .A2(new_n405_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n653_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n539_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n359_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n411_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT122), .B(new_n885_), .C1(new_n827_), .C2(new_n832_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n833_), .A2(KEYINPUT124), .A3(new_n884_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT124), .B1(new_n833_), .B2(new_n884_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n895_), .A2(new_n407_), .A3(new_n714_), .A4(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n886_), .A2(new_n887_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(G169gat), .A3(new_n890_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT123), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n900_), .B2(KEYINPUT62), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n894_), .B2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(KEYINPUT62), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n892_), .A2(new_n893_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n897_), .A4(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n907_), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n867_), .A2(new_n539_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n308_), .A2(G176gat), .A3(new_n883_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n895_), .A2(new_n896_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n308_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n911_), .B1(new_n914_), .B2(new_n410_), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n615_), .A2(new_n450_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT126), .B1(new_n912_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n883_), .A2(new_n616_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n909_), .A2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(G183gat), .B2(new_n920_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n912_), .A2(KEYINPUT126), .A3(new_n917_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n912_), .B2(new_n592_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n824_), .A2(new_n426_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n912_), .B2(new_n925_), .ZN(G1351gat));
  NOR3_X1   g725(.A1(new_n882_), .A2(new_n702_), .A3(new_n539_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n867_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n359_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n431_), .ZN(G1352gat));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n719_), .ZN(new_n931_));
  AND2_X1   g730(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n933_), .ZN(G1353gat));
  INV_X1    g734(.A(new_n928_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n616_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  AND2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  OR3_X1    g740(.A1(new_n928_), .A2(G218gat), .A3(new_n625_), .ZN(new_n942_));
  OAI21_X1  g741(.A(G218gat), .B1(new_n928_), .B2(new_n592_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1355gat));
endmodule


