//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(KEYINPUT77), .A3(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n202_), .B2(KEYINPUT77), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT25), .B1(new_n212_), .B2(KEYINPUT76), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n215_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n207_), .A2(new_n214_), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT77), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n203_), .ZN(new_n224_));
  OR2_X1    g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(KEYINPUT77), .A2(KEYINPUT23), .A3(G183gat), .A4(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n231_), .A3(new_n219_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n222_), .A2(KEYINPUT30), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT30), .B1(new_n222_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT80), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G71gat), .B(G99gat), .Z(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT78), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G227gat), .A3(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G15gat), .B(G43gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT79), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n246_), .B(KEYINPUT79), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n244_), .A3(new_n243_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n228_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n202_), .A2(KEYINPUT77), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n254_));
  INV_X1    g053(.A(new_n215_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n204_), .A4(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n233_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT30), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n222_), .A2(KEYINPUT30), .A3(new_n233_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n236_), .A2(new_n251_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n248_), .A2(new_n250_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n265_), .B(KEYINPUT80), .C1(new_n235_), .C2(new_n234_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268_));
  INV_X1    g067(.A(G134gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G127gat), .ZN(new_n270_));
  INV_X1    g069(.A(G127gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G134gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n272_), .A3(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(G113gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  OAI21_X1  g077(.A(G113gat), .B1(new_n278_), .B2(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n279_), .A3(G120gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(G120gat), .B1(new_n277_), .B2(new_n279_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT31), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n279_), .ZN(new_n285_));
  INV_X1    g084(.A(G120gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n287_), .B2(new_n280_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n267_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n283_), .A2(new_n288_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(KEYINPUT82), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT82), .B1(new_n290_), .B2(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT3), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT2), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n305_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n303_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n299_), .A2(new_n300_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n296_), .B1(new_n311_), .B2(KEYINPUT1), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n299_), .A2(new_n313_), .A3(new_n300_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT29), .B1(new_n307_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT84), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G197gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(G204gat), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322_));
  INV_X1    g121(.A(G204gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(G197gat), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT21), .B1(new_n321_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n324_), .A2(G197gat), .A3(new_n325_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT86), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT21), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT86), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n324_), .A2(new_n333_), .A3(G197gat), .A4(new_n325_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n318_), .A2(new_n320_), .A3(G204gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n331_), .A2(new_n332_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT84), .B(G197gat), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n330_), .A2(KEYINPUT86), .B1(new_n339_), .B2(G204gat), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT87), .A3(new_n332_), .A4(new_n334_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n329_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n334_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n328_), .A2(new_n332_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n316_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n347_), .B(new_n316_), .C1(new_n342_), .C2(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n354_));
  INV_X1    g153(.A(new_n352_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n349_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n312_), .A2(new_n314_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n304_), .A2(new_n306_), .ZN(new_n359_));
  OAI22_X1  g158(.A1(new_n358_), .A2(new_n310_), .B1(new_n359_), .B2(new_n302_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n361_));
  XOR2_X1   g160(.A(G22gat), .B(G50gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT28), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n361_), .B(new_n363_), .Z(new_n364_));
  NAND4_X1  g163(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT88), .A4(new_n355_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n357_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n361_), .B(new_n363_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n353_), .A2(new_n356_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n353_), .A2(KEYINPUT89), .A3(new_n356_), .A4(new_n368_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n295_), .A2(new_n367_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT90), .Z(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT19), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n338_), .A2(new_n341_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n329_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n345_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n258_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n383_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n389_));
  INV_X1    g188(.A(new_n386_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT22), .B(G169gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n392_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n219_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n207_), .A2(new_n225_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n228_), .B(KEYINPUT92), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(KEYINPUT25), .B(G183gat), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n208_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(new_n224_), .A3(new_n226_), .A4(new_n221_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n388_), .A2(new_n389_), .B1(new_n390_), .B2(new_n403_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n342_), .A2(new_n345_), .A3(new_n258_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT91), .B1(new_n405_), .B2(new_n383_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n382_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT94), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT94), .B(new_n258_), .C1(new_n342_), .C2(new_n345_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n403_), .ZN(new_n412_));
  AOI211_X1 g211(.A(new_n383_), .B(new_n381_), .C1(new_n386_), .C2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n378_), .B1(new_n407_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT0), .ZN(new_n418_));
  INV_X1    g217(.A(G57gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G85gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n360_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n307_), .A2(new_n315_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n287_), .A2(new_n424_), .A3(new_n280_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT4), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n360_), .B(new_n427_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n422_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n422_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n421_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT33), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n426_), .A2(new_n428_), .A3(new_n422_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n423_), .A2(new_n425_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n421_), .B1(new_n436_), .B2(new_n430_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n432_), .A2(new_n433_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n384_), .A2(new_n385_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n345_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n387_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n389_), .A3(KEYINPUT20), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n390_), .A2(new_n403_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n406_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n381_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n378_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n414_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n416_), .A2(new_n434_), .A3(new_n438_), .A4(new_n447_), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n429_), .A2(new_n421_), .A3(new_n431_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n432_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n446_), .A2(KEYINPUT32), .ZN(new_n451_));
  AND4_X1   g250(.A1(new_n382_), .A2(new_n406_), .A3(new_n443_), .A4(new_n442_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n398_), .A2(new_n453_), .A3(new_n402_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n383_), .B1(new_n456_), .B2(new_n386_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n382_), .B1(new_n411_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n445_), .A2(new_n414_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n451_), .B(KEYINPUT96), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n450_), .B(new_n459_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n373_), .B1(new_n448_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n367_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n295_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n290_), .A2(new_n292_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n367_), .A2(new_n371_), .A3(new_n372_), .A4(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n450_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT27), .B1(new_n416_), .B2(new_n447_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT98), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n470_), .B(new_n378_), .C1(new_n452_), .C2(new_n458_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n471_), .A2(KEYINPUT27), .A3(new_n447_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n378_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT98), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n469_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n463_), .B1(new_n468_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT72), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT72), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n482_), .B(KEYINPUT14), .C1(new_n478_), .C2(new_n479_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G8gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n487_), .B(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT74), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(KEYINPUT74), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n490_), .B(KEYINPUT15), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n487_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n490_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n498_), .B(new_n493_), .C1(new_n499_), .C2(new_n487_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(G169gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n317_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n477_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n496_), .A2(KEYINPUT75), .A3(new_n500_), .A4(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G230gat), .A2(G233gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT6), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  OR3_X1    g315(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT8), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT10), .B(G99gat), .Z(new_n524_));
  INV_X1    g323(.A(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT64), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(KEYINPUT9), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .A4(new_n515_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(G57gat), .B(G64gat), .Z(new_n535_));
  INV_X1    g334(.A(KEYINPUT11), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n534_), .A3(KEYINPUT11), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT65), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n541_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT65), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n533_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT67), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n523_), .A2(new_n532_), .A3(new_n543_), .A4(new_n546_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT66), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n513_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n533_), .A2(KEYINPUT12), .A3(new_n542_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(new_n512_), .A3(new_n555_), .A4(new_n550_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G120gat), .B(G148gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT68), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT5), .B(G176gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NAND3_X1  g360(.A1(new_n552_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n563_), .A2(new_n564_), .B1(new_n568_), .B2(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n487_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n544_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n212_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G211gat), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n572_), .B2(new_n542_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n579_), .B(KEYINPUT17), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n547_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n572_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n533_), .A2(new_n497_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n523_), .A2(new_n532_), .A3(new_n490_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(KEYINPUT35), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n589_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n595_), .B(new_n594_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT70), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G190gat), .ZN(new_n602_));
  INV_X1    g401(.A(G218gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT71), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n609_), .B2(new_n605_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n605_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n608_), .A3(KEYINPUT71), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n606_), .B1(new_n599_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT37), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n611_), .B(new_n608_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n570_), .A2(new_n587_), .A3(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT73), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT73), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n476_), .B(new_n511_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  AOI21_X1  g424(.A(G1gat), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n450_), .A3(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n624_), .A2(new_n625_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  NAND2_X1  g428(.A1(new_n570_), .A2(new_n510_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n586_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT100), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n606_), .A2(new_n617_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n476_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT101), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n478_), .B1(new_n637_), .B2(new_n450_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n629_), .A2(new_n638_), .A3(KEYINPUT102), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT102), .B1(new_n629_), .B2(new_n638_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1324gat));
  AND2_X1   g440(.A1(new_n416_), .A2(new_n447_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n474_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n471_), .A2(KEYINPUT27), .A3(new_n447_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n642_), .A2(KEYINPUT27), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n623_), .A2(new_n479_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n479_), .B1(new_n637_), .B2(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n646_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n293_), .A2(new_n294_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n623_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n637_), .B2(new_n657_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT103), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(new_n658_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n464_), .B(KEYINPUT104), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n637_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT42), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n623_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n630_), .A2(new_n587_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n476_), .A2(new_n633_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n450_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n448_), .A2(new_n462_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n464_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n295_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n450_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n357_), .A2(new_n366_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n657_), .B1(new_n682_), .B2(new_n372_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n467_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n685_), .B2(new_n645_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(new_n619_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n686_), .A2(KEYINPUT105), .A3(new_n687_), .A4(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n619_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT44), .B1(new_n694_), .B2(new_n674_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(G29gat), .A3(new_n450_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n476_), .A2(KEYINPUT43), .A3(new_n619_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n698_), .B2(KEYINPUT105), .ZN(new_n699_));
  INV_X1    g498(.A(new_n692_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n674_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n694_), .A2(KEYINPUT106), .A3(KEYINPUT44), .A4(new_n674_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n677_), .B1(new_n697_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(G36gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n676_), .A2(new_n707_), .A3(new_n645_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n475_), .B(new_n695_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(new_n707_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT46), .Z(G1329gat));
  INV_X1    g511(.A(new_n705_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n696_), .A2(G43gat), .A3(new_n466_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n676_), .A2(new_n657_), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n713_), .A2(new_n714_), .B1(G43gat), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g516(.A(G50gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n676_), .A2(new_n718_), .A3(new_n669_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n695_), .A2(new_n679_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n705_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n721_), .B2(G50gat), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  AOI211_X1 g522(.A(new_n723_), .B(new_n718_), .C1(new_n705_), .C2(new_n720_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT108), .B(new_n719_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1331gat));
  INV_X1    g528(.A(new_n570_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n510_), .A2(new_n586_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(new_n476_), .A3(new_n688_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n681_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G57gat), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n636_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n681_), .A2(new_n419_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT110), .Z(G1332gat));
  INV_X1    g540(.A(G64gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n738_), .B2(new_n645_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT48), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n742_), .A3(new_n645_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n738_), .B2(new_n657_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n747_), .A3(new_n657_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n738_), .B2(new_n669_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n733_), .A2(new_n753_), .A3(new_n669_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n570_), .A2(new_n587_), .A3(new_n510_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n694_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n681_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n675_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n681_), .A2(G85gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n759_), .B2(new_n475_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n475_), .A2(G92gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  NAND3_X1  g565(.A1(new_n694_), .A2(new_n657_), .A3(new_n758_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n466_), .A2(new_n524_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n767_), .A2(G99gat), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g570(.A1(new_n694_), .A2(new_n464_), .A3(new_n758_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G106gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT52), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n525_), .A3(new_n464_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT112), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n773_), .A2(KEYINPUT52), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n773_), .A2(KEYINPUT52), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n778_), .B(new_n775_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(KEYINPUT53), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(new_n781_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n778_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n645_), .A2(new_n681_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n555_), .A2(new_n550_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT12), .B1(new_n533_), .B2(new_n547_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n513_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n556_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n556_), .A2(new_n792_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n556_), .A2(KEYINPUT114), .A3(new_n792_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n561_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  INV_X1    g599(.A(new_n561_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n556_), .A2(KEYINPUT114), .A3(new_n792_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT114), .B1(new_n556_), .B2(new_n792_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n800_), .B(new_n801_), .C1(new_n804_), .C2(new_n793_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n492_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT115), .B1(new_n806_), .B2(new_n505_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n494_), .B1(new_n487_), .B2(new_n499_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n497_), .B2(new_n487_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(KEYINPUT115), .A3(new_n505_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n810_), .A2(new_n811_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n799_), .A2(new_n805_), .A3(new_n562_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n688_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(KEYINPUT116), .A3(new_n688_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n799_), .A2(new_n805_), .A3(new_n562_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(KEYINPUT58), .A4(new_n812_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT117), .B1(new_n813_), .B2(new_n814_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n818_), .A2(new_n819_), .A3(new_n822_), .A4(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n799_), .A2(new_n805_), .A3(new_n510_), .A4(new_n562_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n812_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n827_), .B2(new_n633_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n829_), .B(new_n634_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n587_), .B1(new_n824_), .B2(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n731_), .A2(KEYINPUT113), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n731_), .A2(KEYINPUT113), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n570_), .A3(new_n619_), .A4(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n684_), .B(new_n788_), .C1(new_n832_), .C2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n822_), .A2(new_n823_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n815_), .B2(new_n688_), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n817_), .B(new_n619_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n828_), .A2(new_n830_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n586_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n836_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n684_), .A4(new_n788_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n839_), .A2(new_n848_), .A3(G113gat), .A4(new_n510_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n276_), .C1(new_n838_), .C2(new_n511_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n846_), .A2(new_n684_), .A3(new_n510_), .A4(new_n788_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n853_), .B2(new_n276_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n849_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT119), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n849_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1340gat));
  INV_X1    g658(.A(new_n838_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n286_), .A2(KEYINPUT60), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n286_), .B1(new_n570_), .B2(KEYINPUT60), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(KEYINPUT120), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n860_), .B(new_n863_), .C1(KEYINPUT120), .C2(new_n862_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n839_), .A2(new_n730_), .A3(new_n848_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n286_), .ZN(G1341gat));
  NOR2_X1   g665(.A1(new_n586_), .A2(new_n271_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n839_), .B(new_n848_), .C1(KEYINPUT121), .C2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G127gat), .B1(new_n868_), .B2(KEYINPUT121), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n587_), .A3(new_n860_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1342gat));
  NAND3_X1  g670(.A1(new_n860_), .A2(new_n269_), .A3(new_n634_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n839_), .A2(new_n688_), .A3(new_n848_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n269_), .ZN(G1343gat));
  NAND3_X1  g673(.A1(new_n846_), .A2(new_n683_), .A3(new_n788_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n511_), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n570_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n586_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT122), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n880_), .B(new_n882_), .ZN(G1346gat));
  OAI21_X1  g682(.A(G162gat), .B1(new_n875_), .B2(new_n619_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n633_), .A2(G162gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n875_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n475_), .A2(new_n450_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n295_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n846_), .A2(new_n668_), .A3(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n511_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT123), .B(new_n887_), .C1(new_n892_), .C2(new_n218_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n218_), .B1(new_n894_), .B2(KEYINPUT62), .ZN(new_n895_));
  OAI221_X1 g694(.A(new_n895_), .B1(new_n894_), .B2(KEYINPUT62), .C1(new_n891_), .C2(new_n511_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n896_), .A3(new_n897_), .ZN(G1348gat));
  OAI21_X1  g697(.A(new_n219_), .B1(new_n891_), .B2(new_n570_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT124), .ZN(new_n900_));
  INV_X1    g699(.A(new_n846_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n464_), .ZN(new_n902_));
  AND4_X1   g701(.A1(G176gat), .A2(new_n902_), .A3(new_n730_), .A4(new_n890_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n900_), .A2(new_n903_), .ZN(G1349gat));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n587_), .A3(new_n890_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n901_), .A2(new_n669_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n889_), .A2(new_n400_), .A3(new_n295_), .A4(new_n586_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n905_), .A2(new_n212_), .B1(new_n906_), .B2(new_n907_), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n891_), .B2(new_n619_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n634_), .A2(new_n208_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT125), .Z(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n891_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1351gat));
  NOR3_X1   g713(.A1(new_n901_), .A2(new_n465_), .A3(new_n889_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n510_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n730_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n324_), .A2(new_n325_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n323_), .B2(new_n918_), .ZN(G1353gat));
  NAND2_X1  g720(.A1(new_n915_), .A2(new_n587_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT63), .B(G211gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n922_), .B2(new_n925_), .ZN(G1354gat));
  NAND2_X1  g725(.A1(new_n915_), .A2(new_n634_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT127), .B(G218gat), .Z(new_n928_));
  NOR2_X1   g727(.A1(new_n619_), .A2(new_n928_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n927_), .A2(new_n928_), .B1(new_n915_), .B2(new_n929_), .ZN(G1355gat));
endmodule


