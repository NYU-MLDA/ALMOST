//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n216_));
  AND4_X1   g015(.A1(new_n206_), .A2(new_n210_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(new_n208_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT64), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n208_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT7), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n218_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n206_), .A3(new_n223_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n213_), .A2(new_n214_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NOR4_X1   g031(.A1(KEYINPUT64), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n225_), .B1(new_n224_), .B2(new_n218_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n203_), .A2(new_n205_), .B1(new_n222_), .B2(KEYINPUT7), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n228_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT8), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G36gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G29gat), .ZN(new_n241_));
  INV_X1    g040(.A(G29gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G36gat), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT70), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT70), .B1(new_n241_), .B2(new_n243_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT71), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT70), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G43gat), .B(G50gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n246_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n246_), .B2(new_n252_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT15), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n253_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT71), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n250_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n246_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT15), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n239_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT72), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n256_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n261_), .A2(KEYINPUT15), .A3(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n239_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n271_));
  NAND2_X1  g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT35), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n261_), .A2(new_n262_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n275_), .B1(new_n239_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(KEYINPUT73), .B(new_n275_), .C1(new_n239_), .C2(new_n276_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n265_), .A2(new_n270_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n273_), .A2(new_n274_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n266_), .A2(new_n267_), .B1(new_n238_), .B2(new_n232_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n284_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G190gat), .B(G218gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G134gat), .B(G162gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n283_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT75), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT77), .ZN(new_n296_));
  INV_X1    g095(.A(new_n282_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n268_), .A2(new_n269_), .A3(new_n239_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n269_), .B1(new_n268_), .B2(new_n239_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n279_), .A2(new_n280_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n297_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT78), .B(new_n296_), .C1(new_n302_), .C2(new_n285_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n285_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n296_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n308_), .A3(new_n291_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n293_), .A2(new_n303_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT37), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT79), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n283_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n305_), .A2(new_n295_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT37), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT37), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G15gat), .B(G22gat), .ZN(new_n322_));
  INV_X1    g121(.A(G1gat), .ZN(new_n323_));
  INV_X1    g122(.A(G8gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT14), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G8gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NAND2_X1  g127(.A1(G231gat), .A2(G233gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(G71gat), .ZN(new_n332_));
  INV_X1    g131(.A(G71gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(KEYINPUT65), .ZN(new_n334_));
  OAI21_X1  g133(.A(G78gat), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(KEYINPUT65), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(G71gat), .ZN(new_n337_));
  INV_X1    g136(.A(G78gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G64gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G57gat), .ZN(new_n341_));
  INV_X1    g140(.A(G57gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G64gat), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n341_), .A2(new_n343_), .A3(KEYINPUT11), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT11), .B1(new_n341_), .B2(new_n343_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n335_), .B(new_n339_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n341_), .A2(new_n343_), .A3(KEYINPUT11), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n338_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n330_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT17), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G127gat), .B(G155gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT16), .ZN(new_n356_));
  XOR2_X1   g155(.A(G183gat), .B(G211gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n354_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n321_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT80), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n206_), .A2(new_n210_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n237_), .B2(KEYINPUT8), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n227_), .A2(KEYINPUT8), .A3(new_n229_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n346_), .A2(new_n350_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n351_), .B1(new_n232_), .B2(new_n238_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n366_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G230gat), .A2(G233gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n370_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n374_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n373_), .A2(KEYINPUT67), .A3(new_n377_), .A4(new_n374_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G120gat), .B(G148gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(G176gat), .B(G204gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .A4(new_n389_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n391_), .A2(KEYINPUT13), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT13), .B1(new_n391_), .B2(new_n392_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n328_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n268_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n261_), .A2(new_n328_), .A3(new_n262_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G229gat), .A2(G233gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n276_), .A2(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n398_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n399_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI211_X1 g204(.A(KEYINPUT81), .B(new_n399_), .C1(new_n402_), .C2(new_n398_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n400_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G113gat), .B(G141gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G169gat), .B(G197gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n400_), .B(new_n410_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n395_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G169gat), .ZN(new_n418_));
  INV_X1    g217(.A(G169gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n420_));
  INV_X1    g219(.A(G176gat), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT83), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT85), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n423_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G183gat), .A2(G190gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT23), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n433_), .B(new_n434_), .C1(G183gat), .C2(G190gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT24), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n427_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT25), .B(G183gat), .ZN(new_n443_));
  INV_X1    g242(.A(G190gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT26), .B1(new_n444_), .B2(KEYINPUT82), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(KEYINPUT26), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n443_), .B(new_n445_), .C1(new_n446_), .C2(KEYINPUT82), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n436_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(G43gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n449_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G127gat), .B(G134gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G120gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n452_), .B(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(G15gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT30), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT31), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n456_), .B(new_n461_), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G218gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G211gat), .ZN(new_n465_));
  INV_X1    g264(.A(G211gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G218gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(G197gat), .B2(G204gat), .ZN(new_n470_));
  INV_X1    g269(.A(G204gat), .ZN(new_n471_));
  INV_X1    g270(.A(G197gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(KEYINPUT89), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n470_), .A3(KEYINPUT21), .A4(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT21), .ZN(new_n475_));
  OAI21_X1  g274(.A(G204gat), .B1(new_n472_), .B2(KEYINPUT89), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n475_), .B(new_n476_), .C1(new_n472_), .C2(G204gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n465_), .A2(new_n467_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(KEYINPUT90), .A2(KEYINPUT21), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n478_), .A2(new_n479_), .B1(KEYINPUT89), .B2(new_n472_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n474_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(G228gat), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G141gat), .ZN(new_n494_));
  INV_X1    g293(.A(G148gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT3), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT3), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(G141gat), .B2(G148gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G141gat), .A2(G148gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n496_), .A2(new_n498_), .B1(new_n500_), .B2(KEYINPUT2), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n490_), .B1(new_n493_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n494_), .A2(new_n495_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n499_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n488_), .B1(KEYINPUT1), .B2(new_n486_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n486_), .A2(KEYINPUT1), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n481_), .B(new_n485_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n485_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n496_), .A2(new_n498_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT2), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n499_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n492_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n500_), .A2(KEYINPUT2), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n491_), .A2(KEYINPUT86), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n512_), .A2(new_n515_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n489_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n507_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n509_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n474_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n511_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n510_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT91), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n510_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n508_), .A2(new_n531_), .A3(new_n509_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n519_), .A2(new_n520_), .A3(new_n509_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT28), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G22gat), .B(G50gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n530_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n538_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT87), .B1(new_n541_), .B2(new_n536_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n537_), .A2(new_n543_), .A3(new_n538_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n529_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n510_), .A2(new_n523_), .A3(KEYINPUT92), .A4(new_n526_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n528_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n540_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G8gat), .B(G36gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G64gat), .B(G92gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G190gat), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n443_), .A2(new_n556_), .B1(new_n441_), .B2(new_n423_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n439_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n438_), .A2(new_n433_), .A3(KEYINPUT93), .A4(new_n434_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT22), .B(G169gat), .Z(new_n562_));
  OAI211_X1 g361(.A(new_n435_), .B(new_n427_), .C1(G176gat), .C2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT20), .B1(new_n564_), .B2(new_n481_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n522_), .B1(new_n436_), .B2(new_n448_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G226gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT19), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n564_), .B2(new_n481_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n436_), .A2(new_n522_), .A3(new_n448_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n570_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n555_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n568_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n561_), .A2(new_n563_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n571_), .B1(new_n578_), .B2(new_n522_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n449_), .A2(new_n481_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n570_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n555_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n577_), .A2(new_n581_), .A3(KEYINPUT95), .A4(new_n582_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n455_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n453_), .B(new_n454_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n519_), .A2(new_n588_), .A3(new_n520_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n589_), .A3(KEYINPUT4), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT4), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n455_), .B(new_n591_), .C1(new_n502_), .C2(new_n507_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(G225gat), .A2(G233gat), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G1gat), .B(G29gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G85gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT0), .B(G57gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n585_), .A2(new_n586_), .B1(new_n595_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n594_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT96), .B1(new_n604_), .B2(new_n600_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT96), .B(KEYINPUT33), .C1(new_n604_), .C2(new_n600_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n582_), .A2(KEYINPUT32), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n577_), .A2(new_n581_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT97), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n604_), .A2(new_n600_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n604_), .A2(new_n600_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n568_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n568_), .B2(new_n576_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(KEYINPUT32), .A3(new_n582_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n550_), .B1(new_n610_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n616_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT27), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n585_), .A2(new_n623_), .A3(new_n586_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n618_), .B2(new_n555_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n583_), .A2(KEYINPUT98), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n577_), .A2(new_n581_), .A3(new_n627_), .A4(new_n582_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  AND4_X1   g428(.A1(new_n550_), .A2(new_n622_), .A3(new_n624_), .A4(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n463_), .B1(new_n621_), .B2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n624_), .A2(new_n629_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n550_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n462_), .A2(new_n632_), .A3(new_n633_), .A4(new_n622_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n416_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n364_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n323_), .A3(new_n616_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n362_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n395_), .A2(new_n415_), .A3(new_n641_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n642_), .A2(KEYINPUT99), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n315_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(KEYINPUT99), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n622_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n638_), .A2(new_n639_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n640_), .A2(new_n647_), .A3(new_n648_), .ZN(G1324gat));
  INV_X1    g448(.A(new_n632_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n637_), .A2(new_n324_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G8gat), .B1(new_n646_), .B2(new_n632_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT100), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(KEYINPUT100), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n651_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT40), .B(new_n651_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n646_), .B2(new_n463_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n637_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT101), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n637_), .A2(new_n668_), .A3(new_n550_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G22gat), .B1(new_n646_), .B2(new_n633_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1327gat));
  OAI21_X1  g471(.A(new_n292_), .B1(new_n305_), .B2(new_n295_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n362_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n636_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n616_), .A2(new_n242_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT105), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n395_), .A2(new_n415_), .A3(new_n362_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT102), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT79), .B1(new_n673_), .B2(KEYINPUT37), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(KEYINPUT37), .B2(new_n310_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT37), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n635_), .B(new_n681_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT104), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n320_), .A2(new_n687_), .A3(new_n681_), .A4(new_n635_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n635_), .A2(new_n690_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n631_), .A2(KEYINPUT103), .A3(new_n634_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n681_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n680_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n680_), .C1(new_n689_), .C2(new_n693_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n696_), .A2(new_n698_), .A3(new_n622_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n678_), .B1(new_n699_), .B2(new_n242_), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n675_), .A2(new_n240_), .A3(new_n650_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT45), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT107), .B1(new_n701_), .B2(KEYINPUT45), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(KEYINPUT107), .A2(G36gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n694_), .A2(new_n695_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n650_), .A3(new_n697_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n706_), .A2(KEYINPUT106), .A3(new_n650_), .A4(new_n697_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT46), .B(new_n704_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n708_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n705_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n710_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n704_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n711_), .A2(new_n717_), .ZN(G1329gat));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n675_), .A2(new_n719_), .A3(new_n462_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n696_), .A2(new_n698_), .A3(new_n463_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n719_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n675_), .B2(new_n550_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n696_), .A2(new_n698_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n550_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(G1331gat));
  INV_X1    g527(.A(new_n395_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n414_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n635_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n364_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n342_), .B1(new_n732_), .B2(new_n622_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT108), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n644_), .A2(new_n362_), .A3(new_n730_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n342_), .A3(new_n622_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n735_), .B2(new_n632_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n650_), .A2(new_n340_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n732_), .B2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n735_), .B2(new_n463_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT49), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n462_), .A2(new_n333_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n732_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n735_), .B2(new_n633_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n550_), .A2(new_n338_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n732_), .B2(new_n748_), .ZN(G1335gat));
  OR2_X1    g548(.A1(new_n689_), .A2(new_n693_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n730_), .A2(new_n641_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n622_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n731_), .A2(new_n674_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n211_), .A3(new_n616_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1336gat));
  OAI21_X1  g557(.A(G92gat), .B1(new_n753_), .B2(new_n632_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n212_), .A3(new_n650_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1337gat));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n207_), .A2(new_n209_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n755_), .A2(new_n763_), .A3(new_n463_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n750_), .A2(new_n462_), .A3(new_n752_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(G99gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n762_), .B1(new_n767_), .B2(KEYINPUT51), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n766_), .A2(KEYINPUT109), .A3(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n766_), .A2(KEYINPUT110), .A3(new_n769_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT110), .B1(new_n766_), .B2(new_n769_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n768_), .A2(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n756_), .A2(new_n208_), .A3(new_n550_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n750_), .A2(new_n550_), .A3(new_n752_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G106gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n650_), .A2(new_n550_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n616_), .A3(new_n462_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n414_), .A2(new_n392_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n232_), .A2(new_n238_), .A3(new_n351_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n365_), .B1(new_n375_), .B2(new_n786_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n239_), .A2(new_n370_), .B1(KEYINPUT66), .B2(KEYINPUT12), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n785_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n373_), .A2(KEYINPUT111), .A3(new_n377_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n381_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n380_), .A2(new_n794_), .A3(new_n383_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n378_), .A2(new_n794_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT112), .A4(new_n381_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n793_), .A2(new_n795_), .A3(new_n796_), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n390_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n390_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n784_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n397_), .A2(new_n398_), .A3(new_n404_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n410_), .B1(new_n403_), .B2(new_n399_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n413_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n673_), .B1(new_n803_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n784_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n390_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n390_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n391_), .A2(new_n392_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n807_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n809_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT113), .B(new_n807_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n315_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT114), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n813_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n819_), .A2(new_n392_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n318_), .A2(new_n319_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT58), .B(new_n827_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n830_), .A2(new_n831_), .B1(new_n823_), .B2(KEYINPUT57), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n362_), .B1(new_n826_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n395_), .A2(new_n414_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(new_n318_), .A3(new_n362_), .A4(new_n319_), .ZN(new_n835_));
  XOR2_X1   g634(.A(new_n835_), .B(KEYINPUT54), .Z(new_n836_));
  OAI21_X1  g635(.A(new_n783_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n414_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n835_), .B(KEYINPUT54), .ZN(new_n841_));
  AOI211_X1 g640(.A(KEYINPUT116), .B(new_n362_), .C1(new_n826_), .C2(new_n832_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n823_), .A2(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n828_), .A2(new_n829_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n320_), .A2(new_n831_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n825_), .B1(new_n823_), .B2(KEYINPUT114), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n812_), .B(new_n315_), .C1(new_n817_), .C2(new_n822_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n844_), .B(new_n846_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n849_), .B2(new_n641_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n841_), .B1(new_n842_), .B2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n782_), .A2(KEYINPUT59), .ZN(new_n852_));
  AOI221_X4 g651(.A(new_n840_), .B1(new_n837_), .B2(KEYINPUT59), .C1(new_n851_), .C2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT117), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n414_), .A2(G113gat), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT118), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n839_), .B1(new_n857_), .B2(new_n859_), .ZN(G1340gat));
  AND3_X1   g659(.A1(new_n854_), .A2(new_n395_), .A3(new_n855_), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(KEYINPUT60), .B2(new_n862_), .ZN(new_n864_));
  OAI22_X1  g663(.A1(new_n861_), .A2(new_n862_), .B1(new_n837_), .B2(new_n864_), .ZN(G1341gat));
  AOI21_X1  g664(.A(G127gat), .B1(new_n838_), .B2(new_n362_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n362_), .A2(G127gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n857_), .B2(new_n867_), .ZN(G1342gat));
  AOI21_X1  g667(.A(G134gat), .B1(new_n838_), .B2(new_n315_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n320_), .A2(G134gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n857_), .B2(new_n870_), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n849_), .A2(new_n641_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n462_), .B1(new_n872_), .B2(new_n841_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(new_n550_), .A3(new_n616_), .A4(new_n632_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n415_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT119), .B(G141gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n875_), .B(new_n876_), .Z(G1344gat));
  NOR2_X1   g676(.A1(new_n874_), .A2(new_n729_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n495_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n874_), .A2(new_n641_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n880_), .B(new_n881_), .Z(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n874_), .B2(new_n321_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n673_), .A2(G162gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n874_), .B2(new_n884_), .ZN(G1347gat));
  NOR3_X1   g684(.A1(new_n463_), .A2(new_n616_), .A3(new_n632_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n550_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n851_), .A2(new_n414_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G169gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n891_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(G169gat), .A3(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n892_), .B(new_n894_), .C1(new_n562_), .C2(new_n889_), .ZN(G1348gat));
  AND2_X1   g694(.A1(new_n851_), .A2(new_n888_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n896_), .B2(new_n395_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n550_), .B1(new_n872_), .B2(new_n841_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n729_), .A2(new_n887_), .A3(new_n421_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n887_), .A2(new_n641_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G183gat), .B1(new_n898_), .B2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n641_), .A2(new_n443_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n896_), .B2(new_n903_), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n896_), .A2(new_n556_), .A3(new_n315_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n851_), .A2(new_n320_), .A3(new_n888_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(G190gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(G190gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n905_), .B1(new_n908_), .B2(new_n909_), .ZN(G1351gat));
  XNOR2_X1  g709(.A(KEYINPUT122), .B(G197gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n472_), .A2(KEYINPUT122), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n650_), .A2(new_n550_), .A3(new_n622_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n873_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n415_), .ZN(new_n916_));
  MUX2_X1   g715(.A(new_n911_), .B(new_n912_), .S(new_n916_), .Z(G1352gat));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n729_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n471_), .A2(KEYINPUT123), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n918_), .B(new_n919_), .Z(G1353gat));
  NOR2_X1   g719(.A1(new_n915_), .A2(new_n641_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT63), .B(G211gat), .Z(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT124), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n921_), .A2(new_n925_), .A3(new_n922_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n915_), .B2(new_n641_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT125), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n930_), .B(new_n927_), .C1(new_n915_), .C2(new_n641_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n924_), .A2(new_n926_), .B1(new_n929_), .B2(new_n931_), .ZN(G1354gat));
  XNOR2_X1  g731(.A(KEYINPUT127), .B(G218gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n915_), .A2(new_n321_), .A3(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n873_), .A2(new_n315_), .A3(new_n914_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT126), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n936_), .B2(new_n933_), .ZN(G1355gat));
endmodule


