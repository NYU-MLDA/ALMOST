//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_;
  NOR3_X1   g000(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n203_), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(KEYINPUT26), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT26), .B(G190gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT77), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT78), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n216_), .B(new_n213_), .C1(new_n221_), .C2(new_n214_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n212_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT80), .B1(new_n208_), .B2(new_n210_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n207_), .B2(KEYINPUT23), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n233_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n225_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n239_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(G15gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n242_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G127gat), .B(G134gat), .Z(new_n249_));
  XOR2_X1   g048(.A(G113gat), .B(G120gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT31), .Z(new_n252_));
  OR2_X1    g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n254_), .A3(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  INV_X1    g057(.A(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT3), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT2), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT82), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(KEYINPUT82), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(KEYINPUT1), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(KEYINPUT1), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n270_), .A2(new_n269_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n263_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n265_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n251_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n272_), .A2(new_n251_), .A3(new_n277_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(KEYINPUT4), .A3(new_n281_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(new_n287_), .A3(new_n279_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n262_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT95), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n262_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n290_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  INV_X1    g099(.A(KEYINPUT94), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT85), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G197gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310_));
  NOR4_X1   g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .A4(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n304_), .A2(new_n306_), .A3(new_n302_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(G197gat), .B2(G204gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT86), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(KEYINPUT86), .A3(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n308_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n310_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT85), .B(G197gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(new_n302_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n322_), .B2(new_n309_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n311_), .B1(new_n318_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n221_), .A2(new_n213_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n206_), .B(new_n325_), .C1(new_n234_), .C2(new_n236_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n211_), .A2(new_n233_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n230_), .B(KEYINPUT93), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n229_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n324_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n311_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n312_), .A2(KEYINPUT86), .A3(new_n313_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT86), .B1(new_n312_), .B2(new_n313_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n304_), .A2(new_n306_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n310_), .B1(new_n337_), .B2(G204gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n308_), .B1(new_n338_), .B2(KEYINPUT21), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n333_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n322_), .A2(new_n309_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(new_n308_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT87), .A3(new_n333_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n222_), .B(new_n223_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n347_), .A2(new_n212_), .B1(new_n237_), .B2(new_n231_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n332_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n301_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  AOI211_X1 g153(.A(new_n341_), .B(new_n311_), .C1(new_n318_), .C2(new_n323_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT87), .B1(new_n344_), .B2(new_n333_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n348_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n332_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT94), .A3(new_n352_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n342_), .A2(new_n239_), .A3(new_n345_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n352_), .B1(new_n324_), .B2(new_n331_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(KEYINPUT20), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n300_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n300_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  AOI211_X1 g166(.A(new_n366_), .B(new_n367_), .C1(new_n354_), .C2(new_n360_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n296_), .B(new_n369_), .C1(new_n295_), .C2(new_n290_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n300_), .A2(KEYINPUT32), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n361_), .A2(new_n371_), .A3(new_n364_), .ZN(new_n372_));
  OR3_X1    g171(.A1(new_n285_), .A2(new_n289_), .A3(new_n262_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n290_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT97), .B1(new_n349_), .B2(new_n353_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n326_), .A2(KEYINPUT96), .A3(new_n329_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT96), .B1(new_n326_), .B2(new_n329_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n340_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n324_), .A2(KEYINPUT89), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n362_), .A3(KEYINPUT20), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n352_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n349_), .A2(new_n353_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n375_), .B1(new_n386_), .B2(KEYINPUT97), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n372_), .B(new_n374_), .C1(new_n387_), .C2(new_n371_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n370_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n390_));
  INV_X1    g189(.A(G233gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT88), .B1(new_n346_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n278_), .B2(KEYINPUT29), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT88), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n342_), .A3(new_n400_), .A4(new_n345_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n380_), .A2(new_n381_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n390_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n395_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n380_), .A2(new_n381_), .B1(KEYINPUT29), .B2(new_n278_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT90), .B1(new_n407_), .B2(new_n396_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n402_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n402_), .A2(new_n406_), .A3(new_n408_), .A4(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G22gat), .B(G50gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  AND4_X1   g217(.A1(KEYINPUT91), .A2(new_n411_), .A3(new_n413_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n421_), .A2(new_n418_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n389_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n374_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT27), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT94), .B1(new_n359_), .B2(new_n352_), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n301_), .B(new_n353_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n300_), .B(new_n364_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT27), .B(new_n431_), .C1(new_n387_), .C2(new_n300_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n423_), .A2(new_n426_), .A3(new_n428_), .A4(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n257_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n428_), .A2(new_n432_), .A3(KEYINPUT98), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT98), .B1(new_n428_), .B2(new_n432_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n424_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT99), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n386_), .A2(KEYINPUT97), .ZN(new_n440_));
  INV_X1    g239(.A(new_n375_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n300_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(KEYINPUT27), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n364_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n366_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT27), .B1(new_n446_), .B2(new_n431_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n439_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n428_), .A2(new_n432_), .A3(KEYINPUT98), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n424_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n438_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n256_), .A2(new_n374_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n434_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT68), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G43gat), .B(G50gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT15), .ZN(new_n460_));
  INV_X1    g259(.A(new_n458_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n457_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT15), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  INV_X1    g264(.A(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n460_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n459_), .A2(new_n471_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n459_), .A2(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G169gat), .B(G197gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n479_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n455_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n496_));
  XOR2_X1   g295(.A(G71gat), .B(G78gat), .Z(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n496_), .A2(new_n497_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(new_n471_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G231gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT73), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n501_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G127gat), .B(G155gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT16), .ZN(new_n507_));
  XOR2_X1   g306(.A(G183gat), .B(G211gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT74), .A3(KEYINPUT17), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n505_), .A2(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n505_), .B(new_n511_), .C1(KEYINPUT17), .C2(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT34), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT35), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n519_), .A2(KEYINPUT70), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n516_), .A2(KEYINPUT35), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G85gat), .B(G92gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT9), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT10), .B(G99gat), .Z(new_n529_));
  INV_X1    g328(.A(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(G85gat), .A3(G92gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT6), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .A4(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  OR3_X1    g335(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n526_), .B1(KEYINPUT65), .B2(KEYINPUT8), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n535_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n525_), .B1(new_n543_), .B2(new_n459_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n547_), .A2(new_n462_), .A3(KEYINPUT69), .A4(new_n535_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n524_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT66), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(KEYINPUT66), .B(new_n535_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n551_), .A2(new_n460_), .A3(new_n464_), .A4(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n522_), .B(new_n523_), .C1(new_n549_), .C2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n549_), .A2(KEYINPUT70), .A3(new_n519_), .A4(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT72), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT71), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n544_), .A2(new_n548_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n524_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n553_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n522_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n523_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n564_), .B1(new_n570_), .B2(new_n555_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n562_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT36), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n555_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n572_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n563_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n563_), .A2(new_n573_), .A3(KEYINPUT37), .A4(new_n575_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n514_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n500_), .B(new_n535_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n500_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n543_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT64), .Z(new_n588_));
  NAND4_X1  g387(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n583_), .A4(new_n552_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n584_), .A2(new_n581_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G120gat), .B(G148gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT5), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n592_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n598_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n580_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n493_), .A2(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n603_), .A2(G1gat), .A3(new_n426_), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n451_), .B1(new_n450_), .B2(new_n424_), .ZN(new_n607_));
  AOI211_X1 g406(.A(KEYINPUT99), .B(new_n423_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n454_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n434_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n576_), .B(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n601_), .A2(new_n491_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n514_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n426_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n604_), .A2(new_n605_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n606_), .A2(new_n618_), .A3(new_n619_), .ZN(G1324gat));
  OAI21_X1  g419(.A(G8gat), .B1(new_n617_), .B2(new_n450_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT39), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n435_), .A2(new_n436_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n493_), .A2(new_n467_), .A3(new_n623_), .A4(new_n602_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g425(.A(G15gat), .B1(new_n617_), .B2(new_n256_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT41), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n603_), .A2(G15gat), .A3(new_n256_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1326gat));
  OAI21_X1  g429(.A(G22gat), .B1(new_n617_), .B2(new_n424_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT42), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n424_), .A2(G22gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n603_), .B2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n514_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n613_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n601_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n493_), .A2(new_n638_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n639_), .A2(G29gat), .A3(new_n426_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n572_), .B1(new_n574_), .B2(KEYINPUT72), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n642_), .A2(new_n558_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT37), .B1(new_n643_), .B2(new_n573_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n579_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n454_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n438_), .B2(new_n452_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n641_), .B(new_n646_), .C1(new_n648_), .C2(new_n434_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n611_), .A2(KEYINPUT102), .A3(new_n641_), .A4(new_n646_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n578_), .A2(new_n579_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n615_), .A2(new_n635_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT44), .B1(new_n655_), .B2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n374_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G29gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n640_), .B1(new_n662_), .B2(new_n663_), .ZN(G1328gat));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n623_), .A2(KEYINPUT104), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n623_), .A2(KEYINPUT104), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n493_), .A2(new_n665_), .A3(new_n638_), .A4(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT45), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n657_), .A2(new_n658_), .A3(new_n450_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n665_), .ZN(new_n672_));
  OR2_X1    g471(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n673_));
  NAND2_X1  g472(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  NAND3_X1  g476(.A1(new_n659_), .A2(G43gat), .A3(new_n257_), .ZN(new_n678_));
  INV_X1    g477(.A(G43gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(new_n639_), .B2(new_n256_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1330gat));
  OR3_X1    g482(.A1(new_n639_), .A2(G50gat), .A3(new_n424_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n659_), .A2(new_n685_), .A3(new_n423_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G50gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n659_), .B2(new_n423_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1331gat));
  NAND4_X1  g488(.A1(new_n614_), .A2(new_n492_), .A3(new_n637_), .A4(new_n635_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n426_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n455_), .A2(new_n491_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n637_), .A3(new_n580_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n426_), .A2(G57gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT108), .ZN(G1332gat));
  INV_X1    g495(.A(new_n668_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G64gat), .B1(new_n690_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT48), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n697_), .A2(G64gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n693_), .B2(new_n700_), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n690_), .B2(new_n256_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n256_), .A2(G71gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n693_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT109), .ZN(G1334gat));
  OAI21_X1  g505(.A(G78gat), .B1(new_n690_), .B2(new_n424_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT50), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n424_), .A2(G78gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n693_), .B2(new_n709_), .ZN(G1335gat));
  NOR3_X1   g509(.A1(new_n601_), .A2(new_n491_), .A3(new_n635_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n655_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n426_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n636_), .A2(new_n601_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n692_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n259_), .A3(new_n374_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1336gat));
  OAI21_X1  g518(.A(G92gat), .B1(new_n713_), .B2(new_n697_), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n716_), .A2(G92gat), .A3(new_n450_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1337gat));
  NAND2_X1  g521(.A1(new_n257_), .A2(new_n529_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n716_), .A2(new_n723_), .B1(KEYINPUT110), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n712_), .A2(new_n257_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G99gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(KEYINPUT110), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n727_), .B(new_n728_), .Z(G1338gat));
  NAND3_X1  g528(.A1(new_n717_), .A2(new_n530_), .A3(new_n423_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n655_), .A2(KEYINPUT111), .A3(new_n423_), .A4(new_n711_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(G106gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n655_), .A2(new_n423_), .A3(new_n711_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n731_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  AND4_X1   g536(.A1(new_n731_), .A2(new_n736_), .A3(G106gat), .A4(new_n732_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n730_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n741_), .B(new_n730_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  NAND2_X1  g542(.A1(new_n602_), .A2(new_n492_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT54), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n590_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n586_), .A2(new_n589_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n588_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n586_), .A2(new_n589_), .A3(KEYINPUT55), .A4(new_n588_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT113), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n596_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n753_), .A2(new_n759_), .A3(KEYINPUT56), .A4(new_n596_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n487_), .B1(new_n481_), .B2(new_n478_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n474_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n490_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n592_), .A2(new_n596_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n761_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n646_), .A2(new_n770_), .A3(KEYINPUT114), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT58), .B1(new_n761_), .B2(new_n767_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n653_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n761_), .A2(KEYINPUT58), .A3(new_n767_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n775_), .A2(new_n776_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n771_), .A2(new_n774_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n758_), .A2(new_n754_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n491_), .C1(new_n592_), .C2(new_n596_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n597_), .A2(new_n490_), .A3(new_n764_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n613_), .A2(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(KEYINPUT116), .A3(new_n786_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n613_), .A2(new_n783_), .A3(KEYINPUT57), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n746_), .B1(new_n792_), .B2(new_n514_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n453_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n794_), .A2(new_n426_), .A3(new_n256_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT59), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT117), .B1(new_n793_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n779_), .A2(new_n786_), .A3(new_n791_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n514_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n746_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT59), .B1(new_n802_), .B2(new_n796_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(new_n791_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n635_), .B1(new_n806_), .B2(new_n790_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n804_), .B(new_n797_), .C1(new_n807_), .C2(new_n746_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n799_), .A2(new_n803_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n492_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n802_), .A2(new_n796_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n492_), .A2(G113gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n810_), .B1(new_n812_), .B2(new_n813_), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n601_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n811_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT118), .ZN(new_n818_));
  OAI21_X1  g617(.A(G120gat), .B1(new_n809_), .B2(new_n601_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n809_), .B2(new_n514_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n514_), .A2(G127gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n812_), .B2(new_n822_), .ZN(G1342gat));
  NAND4_X1  g622(.A1(new_n799_), .A2(new_n646_), .A3(new_n803_), .A4(new_n808_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G134gat), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n812_), .A2(G134gat), .A3(new_n613_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(KEYINPUT119), .A3(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1343gat));
  NOR2_X1   g630(.A1(new_n802_), .A2(new_n257_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n668_), .A2(new_n426_), .A3(new_n424_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n492_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT120), .B(G141gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1344gat));
  NOR2_X1   g636(.A1(new_n834_), .A2(new_n601_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g638(.A1(new_n834_), .A2(new_n514_), .ZN(new_n840_));
  XOR2_X1   g639(.A(KEYINPUT61), .B(G155gat), .Z(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1346gat));
  OAI21_X1  g641(.A(G162gat), .B1(new_n834_), .B2(new_n653_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n613_), .A2(G162gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n834_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT121), .ZN(G1347gat));
  NAND2_X1  g646(.A1(new_n668_), .A2(new_n454_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT122), .Z(new_n849_));
  OAI211_X1 g648(.A(new_n424_), .B(new_n849_), .C1(new_n807_), .C2(new_n746_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n491_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(G169gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n852_), .B2(G169gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n491_), .A2(new_n226_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT123), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n854_), .A2(new_n855_), .B1(new_n850_), .B2(new_n857_), .ZN(G1348gat));
  NOR2_X1   g657(.A1(new_n802_), .A2(new_n423_), .ZN(new_n859_));
  AND4_X1   g658(.A1(G176gat), .A2(new_n859_), .A3(new_n637_), .A4(new_n849_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n227_), .A2(new_n228_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n851_), .B2(new_n637_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n864_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  NOR3_X1   g666(.A1(new_n850_), .A2(new_n213_), .A3(new_n514_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n849_), .A2(new_n635_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G183gat), .B1(new_n859_), .B2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1350gat));
  OR3_X1    g670(.A1(new_n850_), .A2(new_n218_), .A3(new_n613_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G190gat), .B1(new_n850_), .B2(new_n653_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(KEYINPUT125), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(KEYINPUT125), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(G1351gat));
  NOR3_X1   g675(.A1(new_n697_), .A2(new_n374_), .A3(new_n424_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n832_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n492_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n303_), .ZN(G1352gat));
  INV_X1    g679(.A(new_n878_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n637_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n302_), .A2(KEYINPUT126), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1353gat));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n885_));
  INV_X1    g684(.A(G211gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n635_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT127), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n881_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n886_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1354gat));
  OAI21_X1  g690(.A(G218gat), .B1(new_n878_), .B2(new_n653_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n613_), .A2(G218gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n878_), .B2(new_n893_), .ZN(G1355gat));
endmodule


