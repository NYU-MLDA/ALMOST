//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n209_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT65), .A3(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n211_), .A2(new_n220_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  XOR2_X1   g026(.A(G85gat), .B(G92gat), .Z(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NOR4_X1   g028(.A1(new_n216_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(new_n218_), .B2(new_n212_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n208_), .A2(new_n210_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT67), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n211_), .A2(new_n220_), .A3(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(KEYINPUT66), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n228_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT8), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n241_), .B2(new_n228_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n229_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT10), .B(G99gat), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n214_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n249_));
  INV_X1    g048(.A(G85gat), .ZN(new_n250_));
  INV_X1    g049(.A(G92gat), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT9), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n248_), .A2(new_n249_), .A3(new_n252_), .A4(new_n225_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G43gat), .B(G50gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(G29gat), .B(G36gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT15), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT71), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT72), .B1(new_n254_), .B2(new_n259_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n253_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n241_), .A2(new_n228_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT68), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT8), .A3(new_n243_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n267_), .B2(new_n229_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n269_));
  INV_X1    g068(.A(new_n259_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n204_), .A2(new_n205_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n263_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n206_), .B1(new_n262_), .B2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G190gat), .B(G218gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT73), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT74), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n206_), .B(KEYINPUT75), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n261_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n273_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n273_), .A2(new_n282_), .A3(new_n285_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n274_), .B(new_n281_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT37), .ZN(new_n290_));
  OR3_X1    g089(.A1(new_n273_), .A2(new_n282_), .A3(new_n285_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n261_), .B(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n271_), .A2(new_n272_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n263_), .A3(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n286_), .A2(new_n291_), .B1(new_n295_), .B2(new_n206_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n277_), .B(KEYINPUT36), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n289_), .B(new_n290_), .C1(new_n296_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT78), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n274_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n297_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n290_), .A4(new_n289_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n289_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n308_), .B2(new_n290_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(KEYINPUT77), .A3(KEYINPUT37), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n305_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(G1gat), .ZN(new_n313_));
  INV_X1    g112(.A(G8gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT14), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G8gat), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G64gat), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT11), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(KEYINPUT11), .ZN(new_n325_));
  XOR2_X1   g124(.A(G71gat), .B(G78gat), .Z(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n325_), .A2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n322_), .B(new_n329_), .Z(new_n330_));
  AND2_X1   g129(.A1(new_n330_), .A2(KEYINPUT79), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G155gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT16), .ZN(new_n333_));
  XOR2_X1   g132(.A(G183gat), .B(G211gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT17), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n331_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n337_), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n330_), .A2(KEYINPUT17), .A3(new_n336_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n342_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n311_), .A2(KEYINPUT81), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n246_), .A2(new_n329_), .A3(new_n253_), .ZN(new_n348_));
  INV_X1    g147(.A(G230gat), .ZN(new_n349_));
  INV_X1    g148(.A(G233gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT12), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n329_), .B1(new_n246_), .B2(new_n253_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT69), .B(KEYINPUT12), .C1(new_n268_), .C2(new_n329_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n348_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n360_), .A2(new_n355_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n351_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G120gat), .B(G148gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT5), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G176gat), .B(G204gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n362_), .A2(new_n367_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT13), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT13), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n311_), .B2(new_n345_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n346_), .A2(new_n347_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n260_), .A2(new_n320_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n270_), .A2(new_n319_), .A3(new_n318_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G229gat), .A2(G233gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n270_), .B(new_n320_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G113gat), .B(G141gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT83), .ZN(new_n387_));
  XOR2_X1   g186(.A(G169gat), .B(G197gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n385_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT23), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(KEYINPUT23), .B2(new_n392_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(G183gat), .B2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G169gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(new_n399_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n404_), .A2(KEYINPUT21), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(KEYINPUT21), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G197gat), .B(G204gat), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n407_), .A3(KEYINPUT21), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT25), .B(G183gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT26), .B(G190gat), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(KEYINPUT84), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT23), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n392_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n394_), .B2(new_n416_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(KEYINPUT84), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT24), .B1(new_n398_), .B2(new_n399_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421_));
  MUX2_X1   g220(.A(new_n420_), .B(KEYINPUT24), .S(new_n421_), .Z(new_n422_));
  NAND4_X1  g221(.A1(new_n415_), .A2(new_n418_), .A3(new_n419_), .A4(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n403_), .A2(new_n411_), .A3(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n413_), .B(KEYINPUT95), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n412_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n396_), .A3(new_n422_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT96), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT96), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n418_), .B1(G183gat), .B2(G190gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n402_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT20), .B(new_n424_), .C1(new_n432_), .C2(new_n411_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT19), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n403_), .A2(new_n423_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n410_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n435_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n411_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n433_), .A2(new_n435_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G8gat), .B(G36gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT98), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n442_), .A2(new_n448_), .ZN(new_n450_));
  MUX2_X1   g249(.A(new_n449_), .B(KEYINPUT98), .S(new_n450_), .Z(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(KEYINPUT27), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT1), .ZN(new_n454_));
  OR2_X1    g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(KEYINPUT1), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(new_n457_), .B2(new_n456_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n454_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n460_), .B2(new_n459_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G141gat), .A2(G148gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT88), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT91), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n466_), .B(KEYINPUT3), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n469_), .B(new_n470_), .C1(new_n465_), .C2(KEYINPUT2), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n455_), .A2(new_n453_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n462_), .A2(new_n467_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G134gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G120gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n473_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(KEYINPUT99), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(new_n476_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n479_), .B2(KEYINPUT4), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT100), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT0), .ZN(new_n487_));
  INV_X1    g286(.A(G57gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n250_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n490_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n483_), .A2(new_n484_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n442_), .A2(new_n448_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n433_), .A2(new_n435_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n410_), .B(KEYINPUT93), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n439_), .B1(new_n498_), .B2(new_n438_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n495_), .B(KEYINPUT27), .C1(new_n500_), .C2(new_n448_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n452_), .A2(new_n494_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n437_), .B(KEYINPUT30), .ZN(new_n504_));
  XOR2_X1   g303(.A(G71gat), .B(G99gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G15gat), .B(G43gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT86), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n507_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n504_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT31), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n476_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT31), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n511_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n476_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT87), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n473_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(G228gat), .B(G233gat), .C1(new_n521_), .C2(new_n497_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n411_), .B1(G228gat), .B2(G233gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n473_), .B2(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G78gat), .B(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n525_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT94), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n473_), .A2(new_n520_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT28), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G22gat), .B(G50gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n530_), .B(new_n534_), .C1(KEYINPUT94), .C2(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(KEYINPUT94), .C1(new_n528_), .C2(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n519_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(new_n518_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n503_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n519_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n493_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n493_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n480_), .A2(new_n481_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n492_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AND4_X1   g348(.A1(new_n451_), .A2(new_n545_), .A3(new_n546_), .A4(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n448_), .A2(KEYINPUT32), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n500_), .A2(KEYINPUT101), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n442_), .B2(new_n551_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT101), .B1(new_n500_), .B2(new_n551_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(new_n494_), .A3(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n543_), .B(new_n538_), .C1(new_n550_), .C2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n542_), .A2(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n377_), .A2(new_n391_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n346_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT82), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n313_), .A3(new_n494_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT38), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n308_), .A2(new_n345_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n375_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n391_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n494_), .ZN(new_n572_));
  OAI21_X1  g371(.A(G1gat), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n563_), .A2(new_n573_), .ZN(G1324gat));
  NOR2_X1   g373(.A1(new_n452_), .A2(new_n502_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(G8gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n558_), .A2(new_n560_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT102), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT102), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n558_), .A2(new_n579_), .A3(new_n560_), .A4(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n575_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n314_), .B1(new_n570_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(KEYINPUT103), .A3(KEYINPUT39), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT103), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n586_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n585_), .B(new_n588_), .C1(KEYINPUT39), .C2(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n581_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT40), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n581_), .A2(new_n589_), .A3(KEYINPUT40), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1325gat));
  INV_X1    g393(.A(G15gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n561_), .A2(new_n595_), .A3(new_n519_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n570_), .B2(new_n519_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT41), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(G1326gat));
  INV_X1    g398(.A(G22gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n561_), .A2(new_n600_), .A3(new_n540_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n570_), .B2(new_n540_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT42), .Z(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(G1327gat));
  INV_X1    g403(.A(new_n345_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n307_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n557_), .A2(new_n568_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(G29gat), .B1(new_n607_), .B2(new_n494_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n557_), .A2(new_n311_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT43), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n557_), .A2(new_n611_), .A3(new_n311_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n605_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(KEYINPUT44), .A3(new_n568_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n614_), .A2(G29gat), .A3(new_n494_), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n569_), .B(new_n605_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n608_), .B1(new_n615_), .B2(new_n620_), .ZN(G1328gat));
  OAI211_X1 g420(.A(new_n614_), .B(new_n582_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G36gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n607_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n624_), .A2(G36gat), .A3(new_n575_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT46), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(KEYINPUT46), .A3(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1329gat));
  INV_X1    g431(.A(new_n518_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(G43gat), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n614_), .B(new_n634_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G43gat), .B1(new_n607_), .B2(new_n519_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT106), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g438(.A1(new_n614_), .A2(G50gat), .A3(new_n540_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n624_), .A2(new_n538_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n640_), .A2(new_n619_), .B1(G50gat), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1331gat));
  NOR3_X1   g443(.A1(new_n565_), .A2(new_n391_), .A3(new_n375_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G57gat), .B1(new_n646_), .B2(new_n572_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n375_), .A2(new_n391_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n557_), .A2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(new_n376_), .A3(new_n346_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n488_), .A3(new_n494_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n651_), .ZN(G1332gat));
  INV_X1    g451(.A(G64gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n645_), .B2(new_n582_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n653_), .A3(new_n582_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g458(.A(G71gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n645_), .B2(new_n519_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT49), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n650_), .A2(new_n660_), .A3(new_n519_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1334gat));
  INV_X1    g463(.A(G78gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n645_), .B2(new_n540_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT50), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n540_), .A2(new_n665_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT110), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n650_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1335gat));
  NAND2_X1  g470(.A1(new_n613_), .A2(new_n648_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n613_), .A2(KEYINPUT111), .A3(new_n648_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n250_), .B1(new_n676_), .B2(new_n494_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n649_), .A2(new_n606_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n494_), .A2(new_n250_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT112), .B1(new_n677_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT112), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n572_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n683_));
  OAI221_X1 g482(.A(new_n682_), .B1(new_n678_), .B2(new_n679_), .C1(new_n683_), .C2(new_n250_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1336gat));
  INV_X1    g484(.A(new_n678_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n251_), .A3(new_n582_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n575_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n251_), .ZN(G1337gat));
  AOI21_X1  g488(.A(new_n213_), .B1(new_n676_), .B2(new_n519_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n633_), .A2(new_n247_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n678_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT51), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT51), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n543_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n695_));
  OAI221_X1 g494(.A(new_n694_), .B1(new_n678_), .B2(new_n691_), .C1(new_n695_), .C2(new_n213_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1338gat));
  NAND3_X1  g496(.A1(new_n686_), .A2(new_n214_), .A3(new_n540_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n613_), .A2(new_n540_), .A3(new_n648_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT52), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(G106gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G106gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(G1339gat));
  NAND2_X1  g504(.A1(new_n575_), .A2(new_n494_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n541_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT59), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n309_), .A2(new_n310_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n305_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT114), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n345_), .A2(new_n391_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n375_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n375_), .B2(new_n716_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n714_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT54), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n390_), .B1(new_n384_), .B2(new_n381_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n380_), .B(KEYINPUT115), .Z(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n381_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n385_), .A2(new_n390_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n369_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n360_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(KEYINPUT55), .A2(new_n359_), .B1(new_n729_), .B2(new_n352_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n359_), .A2(KEYINPUT55), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n366_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT56), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT118), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT56), .B(new_n366_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n729_), .A2(new_n352_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n359_), .A2(KEYINPUT55), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n359_), .A2(KEYINPUT55), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n366_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT118), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n728_), .B1(new_n737_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT119), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT58), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n735_), .B1(new_n742_), .B2(KEYINPUT118), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n732_), .A2(KEYINPUT118), .A3(new_n733_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n727_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(KEYINPUT119), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n746_), .A2(new_n311_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n368_), .A2(new_n391_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n732_), .A2(new_n733_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n735_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n726_), .B1(new_n372_), .B2(new_n368_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n307_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n753_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n742_), .B2(new_n736_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n756_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n308_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT57), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n752_), .A2(new_n759_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n345_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n711_), .B1(new_n721_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n759_), .A2(new_n768_), .B1(KEYINPUT57), .B2(new_n763_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n757_), .A2(KEYINPUT117), .A3(new_n758_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n752_), .A2(KEYINPUT120), .A3(new_n769_), .A4(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n345_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n758_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n763_), .B2(new_n773_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n774_), .A2(new_n770_), .A3(new_n764_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT120), .B1(new_n775_), .B2(new_n752_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n721_), .B1(new_n772_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n709_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n767_), .B1(new_n778_), .B2(KEYINPUT59), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G113gat), .B1(new_n780_), .B2(new_n567_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n567_), .A2(G113gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n778_), .B2(new_n782_), .ZN(G1340gat));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT121), .B(G120gat), .Z(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n779_), .B2(new_n566_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT60), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n566_), .A2(new_n787_), .A3(new_n785_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT60), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n778_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n767_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n775_), .A2(new_n752_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n345_), .A3(new_n771_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n708_), .B1(new_n797_), .B2(new_n721_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n566_), .B(new_n793_), .C1(new_n798_), .C2(new_n710_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n789_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n791_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(KEYINPUT122), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n792_), .A2(new_n802_), .ZN(G1341gat));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n804_));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n779_), .B2(new_n605_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n778_), .A2(G127gat), .A3(new_n345_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n804_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n605_), .B(new_n793_), .C1(new_n798_), .C2(new_n710_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G127gat), .ZN(new_n810_));
  INV_X1    g609(.A(new_n807_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(KEYINPUT123), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n812_), .ZN(G1342gat));
  OAI21_X1  g612(.A(G134gat), .B1(new_n780_), .B2(new_n714_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n307_), .A2(G134gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n778_), .B2(new_n815_), .ZN(G1343gat));
  AND2_X1   g615(.A1(new_n777_), .A2(new_n539_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n391_), .A3(new_n707_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n566_), .A3(new_n707_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n707_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n345_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT61), .B(G155gat), .Z(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  OAI21_X1  g624(.A(G162gat), .B1(new_n822_), .B2(new_n714_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n307_), .A2(G162gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n822_), .B2(new_n827_), .ZN(G1347gat));
  NAND2_X1  g627(.A1(new_n721_), .A2(new_n766_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n575_), .A2(new_n494_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n519_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n540_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n391_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G169gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n829_), .A2(new_n832_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n391_), .A3(new_n401_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n836_), .A2(new_n839_), .A3(KEYINPUT124), .A4(new_n837_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1348gat));
  AOI21_X1  g643(.A(G176gat), .B1(new_n838_), .B2(new_n566_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(KEYINPUT125), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(KEYINPUT125), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n540_), .B1(new_n797_), .B2(new_n721_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n831_), .A2(new_n399_), .A3(new_n375_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n846_), .A2(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(G1349gat));
  NAND4_X1  g649(.A1(new_n848_), .A2(new_n519_), .A3(new_n605_), .A4(new_n830_), .ZN(new_n851_));
  INV_X1    g650(.A(G183gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n345_), .A2(new_n412_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n851_), .A2(new_n852_), .B1(new_n838_), .B2(new_n853_), .ZN(G1350gat));
  NAND2_X1  g653(.A1(new_n838_), .A2(new_n311_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G190gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n838_), .A2(new_n425_), .A3(new_n308_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1351gat));
  NAND2_X1  g657(.A1(new_n817_), .A2(new_n830_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n567_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT126), .B(G197gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1352gat));
  INV_X1    g661(.A(G204gat), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n863_), .A2(KEYINPUT127), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n817_), .A2(new_n566_), .A3(new_n830_), .A4(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(KEYINPUT127), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1353gat));
  NOR2_X1   g666(.A1(new_n859_), .A2(new_n345_), .ZN(new_n868_));
  AND2_X1   g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n868_), .B2(new_n870_), .ZN(G1354gat));
  OAI21_X1  g672(.A(G218gat), .B1(new_n859_), .B2(new_n714_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n307_), .A2(G218gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n859_), .B2(new_n875_), .ZN(G1355gat));
endmodule


