//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n989_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT82), .B(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT22), .B(G169gat), .ZN(new_n213_));
  AOI211_X1 g012(.A(KEYINPUT83), .B(new_n211_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT82), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G169gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n217_), .A2(new_n219_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n215_), .B1(new_n224_), .B2(new_n210_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n209_), .B1(new_n214_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n220_), .A2(new_n216_), .A3(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT24), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n204_), .A2(new_n208_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n227_), .A2(new_n229_), .A3(KEYINPUT24), .A4(new_n210_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n206_), .A2(KEYINPUT26), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G190gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT80), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT25), .B(G183gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(KEYINPUT80), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n232_), .B(new_n233_), .C1(new_n237_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n226_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G15gat), .B(G43gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G134gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G127gat), .ZN(new_n255_));
  INV_X1    g054(.A(G127gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G134gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n253_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n256_), .A2(G134gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n254_), .A2(G127gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT85), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n252_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT31), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n251_), .B1(KEYINPUT86), .B2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n243_), .A2(new_n244_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n269_), .B(new_n271_), .C1(KEYINPUT86), .C2(new_n268_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  INV_X1    g072(.A(new_n268_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n271_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(new_n274_), .C1(new_n275_), .C2(new_n251_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT91), .ZN(new_n277_));
  INV_X1    g076(.A(G197gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(G204gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(G204gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT21), .ZN(new_n284_));
  INV_X1    g083(.A(G218gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G211gat), .ZN(new_n286_));
  INV_X1    g085(.A(G211gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G218gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n284_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT92), .B1(new_n283_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n283_), .A2(new_n289_), .A3(KEYINPUT92), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n286_), .A2(new_n288_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n281_), .A2(G197gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n280_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(KEYINPUT21), .B2(new_n296_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n291_), .A2(new_n292_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299_));
  OR2_X1    g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(new_n300_), .B2(KEYINPUT87), .ZN(new_n301_));
  NOR3_X1   g100(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT2), .B1(new_n305_), .B2(KEYINPUT88), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n301_), .A2(new_n304_), .A3(new_n306_), .A4(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311_));
  AND2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G155gat), .ZN(new_n315_));
  INV_X1    g114(.A(G162gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(KEYINPUT89), .A3(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n300_), .B(new_n322_), .C1(new_n323_), .C2(new_n318_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT1), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n299_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(G228gat), .B(G233gat), .C1(new_n298_), .C2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n297_), .B1(KEYINPUT21), .B2(new_n283_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n292_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(new_n331_), .B2(new_n290_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n326_), .B1(new_n310_), .B2(new_n320_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n332_), .B(new_n333_), .C1(new_n334_), .C2(new_n299_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  NAND2_X1  g135(.A1(new_n321_), .A2(new_n327_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(KEYINPUT29), .ZN(new_n338_));
  INV_X1    g137(.A(new_n336_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n299_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n329_), .B(new_n335_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n329_), .A2(new_n335_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n344_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n314_), .A2(new_n319_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n302_), .B(KEYINPUT3), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n307_), .B(KEYINPUT2), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n267_), .B1(new_n357_), .B2(new_n326_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n321_), .A2(new_n327_), .A3(new_n266_), .A4(new_n261_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n337_), .A2(new_n363_), .A3(new_n267_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n358_), .A2(new_n361_), .A3(new_n359_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n368_));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n362_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n372_), .B(new_n366_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n272_), .A2(new_n276_), .A3(new_n353_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n227_), .A2(new_n229_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n384_));
  INV_X1    g183(.A(new_n231_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n205_), .A2(KEYINPUT25), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G183gat), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n234_), .A2(new_n236_), .A3(new_n387_), .A4(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n233_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT93), .B1(new_n230_), .B2(new_n231_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n386_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n209_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n204_), .A2(new_n207_), .A3(KEYINPUT94), .A4(new_n208_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n332_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n298_), .A2(new_n226_), .A3(new_n241_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .A4(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n399_), .B2(new_n332_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n209_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n224_), .A2(new_n210_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT83), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n394_), .A2(new_n215_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n407_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n233_), .B1(new_n240_), .B2(new_n237_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n383_), .A2(new_n385_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n332_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT95), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n332_), .B(new_n417_), .C1(new_n411_), .C2(new_n414_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n406_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n405_), .B1(new_n419_), .B2(new_n404_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT18), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G64gat), .ZN(new_n423_));
  INV_X1    g222(.A(G92gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n420_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT99), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n429_));
  INV_X1    g228(.A(new_n398_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n233_), .A2(new_n390_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n413_), .B2(KEYINPUT93), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n432_), .B2(new_n386_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n433_), .B2(new_n298_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n418_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n417_), .B1(new_n242_), .B2(new_n332_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n434_), .B(new_n404_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n403_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n425_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT99), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n420_), .A2(new_n441_), .A3(new_n426_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n428_), .A2(KEYINPUT27), .A3(new_n440_), .A4(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n437_), .A2(new_n425_), .A3(new_n439_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n425_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n380_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n437_), .A2(new_n439_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n426_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n377_), .A2(KEYINPUT33), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n365_), .A2(new_n453_), .A3(new_n372_), .A4(new_n366_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n364_), .A2(new_n361_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n372_), .B1(new_n456_), .B2(new_n360_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n358_), .A2(KEYINPUT97), .A3(new_n359_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT97), .B1(new_n358_), .B2(new_n359_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n362_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n451_), .A2(new_n455_), .A3(new_n440_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT98), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n452_), .A2(new_n454_), .B1(new_n460_), .B2(new_n457_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n440_), .A4(new_n451_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n420_), .A2(new_n468_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n463_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n353_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT100), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n352_), .A2(new_n379_), .A3(new_n447_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n420_), .A2(new_n441_), .A3(new_n426_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n441_), .B1(new_n420_), .B2(new_n426_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n440_), .A2(KEYINPUT27), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n474_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n350_), .A2(new_n351_), .A3(new_n378_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n443_), .A2(KEYINPUT100), .A3(new_n481_), .A4(new_n447_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n272_), .A2(new_n276_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n449_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n486_));
  INV_X1    g285(.A(G230gat), .ZN(new_n487_));
  INV_X1    g286(.A(G233gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n494_), .A2(new_n497_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT8), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n504_), .A3(new_n501_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n506_));
  INV_X1    g305(.A(G85gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT64), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT64), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G85gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n424_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n506_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n516_), .A3(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n497_), .A2(new_n498_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n503_), .A2(new_n505_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT11), .ZN(new_n521_));
  INV_X1    g320(.A(G57gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(G64gat), .ZN(new_n523_));
  INV_X1    g322(.A(G64gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(G57gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(G57gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n522_), .A2(G64gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(KEYINPUT11), .ZN(new_n529_));
  XOR2_X1   g328(.A(G71gat), .B(G78gat), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G71gat), .B(G78gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n532_), .A2(KEYINPUT11), .A3(new_n527_), .A4(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n490_), .B1(new_n520_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n514_), .A2(new_n519_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n500_), .A2(new_n504_), .A3(new_n501_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n504_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n534_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(KEYINPUT66), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n534_), .B(new_n536_), .C1(new_n538_), .C2(new_n537_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT65), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n503_), .A2(new_n505_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n546_), .A2(KEYINPUT65), .A3(new_n534_), .A4(new_n536_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n489_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n520_), .A2(new_n534_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n550_), .A2(new_n551_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n539_), .B(new_n540_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n489_), .B1(new_n520_), .B2(new_n534_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n281_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT5), .B(G176gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  AND3_X1   g360(.A1(new_n549_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n549_), .B2(new_n557_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n561_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n489_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n520_), .A2(new_n490_), .A3(new_n534_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT66), .B1(new_n539_), .B2(new_n540_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n545_), .A2(new_n547_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n567_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n557_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n566_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n549_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT68), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n486_), .B1(new_n565_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n564_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(KEYINPUT68), .A3(new_n575_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT13), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT77), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  XNOR2_X1  g389(.A(G29gat), .B(G36gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G43gat), .B(G50gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G29gat), .B(G36gat), .Z(new_n594_));
  XOR2_X1   g393(.A(G43gat), .B(G50gat), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G1gat), .A2(G8gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT14), .ZN(new_n598_));
  NOR2_X1   g397(.A1(G15gat), .A2(G22gat), .ZN(new_n599_));
  AND2_X1   g398(.A1(G15gat), .A2(G22gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(G1gat), .ZN(new_n602_));
  INV_X1    g401(.A(G8gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n597_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G15gat), .B(G22gat), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n607_), .A2(new_n598_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n593_), .B(new_n596_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n601_), .A2(new_n605_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n607_), .A2(new_n597_), .A3(new_n604_), .A4(new_n598_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n593_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n591_), .A2(new_n592_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n610_), .B(new_n611_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(new_n614_), .A3(KEYINPUT76), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n596_), .A2(new_n593_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n610_), .A2(new_n611_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT76), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n615_), .A2(new_n617_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT15), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n596_), .A2(KEYINPUT15), .A3(new_n593_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n620_), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n616_), .A3(new_n614_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n590_), .B1(new_n623_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n628_), .A3(new_n590_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(KEYINPUT78), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(KEYINPUT78), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(KEYINPUT78), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT79), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n631_), .A2(KEYINPUT78), .A3(new_n632_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n629_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n485_), .A2(new_n586_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT37), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n539_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT70), .Z(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT34), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT35), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n643_), .B(new_n648_), .C1(new_n539_), .C2(new_n619_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT36), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n654_), .B(KEYINPUT36), .Z(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n651_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT71), .B(new_n642_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n642_), .A2(KEYINPUT71), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n642_), .A2(KEYINPUT71), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n662_), .A2(new_n656_), .A3(new_n663_), .A4(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n606_), .A2(new_n608_), .A3(KEYINPUT72), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT72), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n669_));
  INV_X1    g468(.A(G231gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n488_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n667_), .A2(new_n669_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT72), .B1(new_n606_), .B2(new_n608_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n610_), .A2(new_n611_), .A3(new_n668_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n534_), .B1(new_n672_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(G183gat), .B(G211gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G127gat), .B(G155gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT17), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n671_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n674_), .A2(new_n675_), .A3(new_n673_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n540_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n677_), .A2(new_n684_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT74), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT74), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n677_), .A2(new_n684_), .A3(new_n687_), .A4(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n682_), .B(KEYINPUT17), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n677_), .A2(new_n687_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT75), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(KEYINPUT75), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n666_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n641_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT101), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT38), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n378_), .A2(new_n602_), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n657_), .A2(new_n660_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n485_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n700_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n640_), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n709_), .A2(new_n584_), .A3(new_n585_), .A4(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G1gat), .B1(new_n712_), .B2(new_n379_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n713_), .A3(new_n714_), .ZN(G1324gat));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n448_), .A3(new_n711_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n603_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n448_), .A2(new_n603_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n721_), .A2(new_n722_), .B1(new_n703_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT40), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI221_X1 g525(.A(KEYINPUT40), .B1(new_n703_), .B2(new_n723_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1325gat));
  OAI21_X1  g527(.A(G15gat), .B1(new_n712_), .B2(new_n484_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT104), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT104), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n703_), .A2(G15gat), .A3(new_n484_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(KEYINPUT41), .A3(new_n731_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(G1326gat));
  OAI21_X1  g536(.A(G22gat), .B1(new_n712_), .B2(new_n353_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT42), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT42), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n353_), .A2(G22gat), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n739_), .A2(new_n740_), .B1(new_n703_), .B2(new_n741_), .ZN(G1327gat));
  AND2_X1   g541(.A1(new_n700_), .A2(new_n707_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n641_), .A2(new_n743_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n744_), .A2(G29gat), .A3(new_n379_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n584_), .A2(new_n700_), .A3(new_n585_), .A4(new_n710_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n480_), .A2(new_n482_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n462_), .A2(KEYINPUT98), .B1(new_n470_), .B2(new_n469_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n352_), .B1(new_n748_), .B2(new_n466_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n484_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n449_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n666_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n666_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n485_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n746_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n378_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n746_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n753_), .B1(new_n752_), .B2(new_n666_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n485_), .A2(KEYINPUT43), .A3(new_n755_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT44), .B(new_n760_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n757_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n759_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768_));
  OAI21_X1  g567(.A(G29gat), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n758_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n770_), .A2(new_n768_), .A3(new_n378_), .A4(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n745_), .B1(new_n769_), .B2(new_n775_), .ZN(G1328gat));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n777_));
  INV_X1    g576(.A(G36gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n448_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n770_), .B2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n448_), .B(KEYINPUT108), .Z(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n778_), .ZN(new_n784_));
  OR3_X1    g583(.A1(new_n744_), .A2(KEYINPUT45), .A3(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT45), .B1(new_n744_), .B2(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n777_), .B1(new_n781_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n779_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT46), .B(new_n787_), .C1(new_n790_), .C2(new_n778_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1329gat));
  XNOR2_X1  g591(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n744_), .A2(new_n484_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n765_), .A2(new_n766_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n484_), .ZN(new_n796_));
  OAI211_X1 g595(.A(G43gat), .B(new_n796_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n797_));
  OAI221_X1 g596(.A(new_n793_), .B1(G43gat), .B2(new_n794_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n793_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n794_), .A2(G43gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(G1330gat));
  INV_X1    g602(.A(new_n744_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G50gat), .B1(new_n804_), .B2(new_n352_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n773_), .A2(G50gat), .A3(new_n352_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n770_), .ZN(G1331gat));
  AND3_X1   g606(.A1(new_n698_), .A2(new_n640_), .A3(new_n699_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n586_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n708_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G57gat), .B1(new_n810_), .B2(new_n379_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n485_), .A2(new_n710_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT110), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n586_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n814_), .A2(new_n700_), .A3(new_n666_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n378_), .A2(new_n522_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n816_), .B2(new_n817_), .ZN(G1332gat));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n524_), .A3(new_n783_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G64gat), .B1(new_n810_), .B2(new_n782_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(KEYINPUT48), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(KEYINPUT48), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n819_), .B1(new_n821_), .B2(new_n822_), .ZN(G1333gat));
  OAI21_X1  g622(.A(G71gat), .B1(new_n810_), .B2(new_n484_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n824_), .A2(KEYINPUT111), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT111), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n825_), .A2(KEYINPUT49), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT49), .B1(new_n825_), .B2(new_n826_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n484_), .A2(G71gat), .ZN(new_n829_));
  OAI22_X1  g628(.A1(new_n827_), .A2(new_n828_), .B1(new_n816_), .B2(new_n829_), .ZN(G1334gat));
  NOR2_X1   g629(.A1(new_n353_), .A2(G78gat), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n813_), .A2(new_n701_), .A3(new_n586_), .A4(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n708_), .A2(new_n809_), .A3(new_n352_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(G78gat), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(new_n833_), .A3(G78gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1335gat));
  NAND3_X1  g638(.A1(new_n586_), .A2(new_n700_), .A3(new_n640_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n379_), .B(new_n842_), .C1(new_n508_), .C2(new_n510_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n813_), .A2(new_n586_), .A3(new_n378_), .A4(new_n743_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n507_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(KEYINPUT113), .A3(new_n507_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n843_), .B1(new_n847_), .B2(new_n848_), .ZN(G1336gat));
  INV_X1    g648(.A(new_n814_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(new_n424_), .A3(new_n448_), .A4(new_n743_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G92gat), .B1(new_n842_), .B2(new_n782_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1337gat));
  NOR2_X1   g652(.A1(new_n842_), .A2(new_n484_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n492_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n484_), .A2(new_n516_), .A3(new_n515_), .ZN(new_n856_));
  AND4_X1   g655(.A1(new_n586_), .A2(new_n813_), .A3(new_n743_), .A4(new_n856_), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n855_), .A2(new_n857_), .A3(KEYINPUT51), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT51), .B1(new_n855_), .B2(new_n857_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1338gat));
  NOR2_X1   g659(.A1(new_n353_), .A2(G106gat), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n813_), .A2(new_n586_), .A3(new_n743_), .A4(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n841_), .A2(new_n352_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(G106gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n863_), .ZN(new_n866_));
  AOI211_X1 g665(.A(new_n493_), .B(new_n866_), .C1(new_n841_), .C2(new_n352_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n862_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT53), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n862_), .C1(new_n865_), .C2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1339gat));
  INV_X1    g671(.A(new_n590_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n615_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n627_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n876_), .A2(new_n631_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n575_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n552_), .A2(new_n555_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n489_), .B1(new_n879_), .B2(new_n548_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n557_), .A2(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .A4(KEYINPUT55), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n884_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n884_), .B2(new_n566_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n878_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT58), .B(new_n878_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n666_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n710_), .B(new_n575_), .C1(new_n886_), .C2(new_n885_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n578_), .A2(new_n579_), .A3(new_n877_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n707_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n891_), .B1(new_n894_), .B2(KEYINPUT57), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n896_), .B(new_n707_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n700_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT13), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT13), .B1(new_n578_), .B2(new_n579_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n808_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n808_), .B(KEYINPUT115), .C1(new_n900_), .C2(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n899_), .B1(new_n906_), .B2(new_n755_), .ZN(new_n907_));
  AOI211_X1 g706(.A(KEYINPUT54), .B(new_n666_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n898_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n448_), .A2(new_n484_), .A3(new_n379_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n353_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(G113gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n913_), .A3(new_n710_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(KEYINPUT59), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n909_), .A2(new_n916_), .A3(new_n353_), .A4(new_n910_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(new_n710_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n914_), .B1(new_n919_), .B2(new_n913_), .ZN(G1340gat));
  NAND3_X1  g719(.A1(new_n915_), .A2(new_n586_), .A3(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(G120gat), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923_));
  INV_X1    g722(.A(new_n586_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(G120gat), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n912_), .B(new_n925_), .C1(new_n923_), .C2(G120gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT116), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT116), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n922_), .A2(new_n929_), .A3(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1341gat));
  NAND3_X1  g730(.A1(new_n912_), .A2(new_n256_), .A3(new_n709_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n918_), .A2(new_n709_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n256_), .ZN(G1342gat));
  AOI21_X1  g733(.A(G134gat), .B1(new_n912_), .B2(new_n707_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n666_), .A2(G134gat), .ZN(new_n936_));
  XOR2_X1   g735(.A(new_n936_), .B(KEYINPUT117), .Z(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n918_), .B2(new_n937_), .ZN(G1343gat));
  NOR2_X1   g737(.A1(new_n796_), .A2(new_n353_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n909_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n783_), .A2(new_n379_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n710_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n586_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT118), .B(G148gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n946_), .B(new_n947_), .ZN(G1345gat));
  INV_X1    g747(.A(new_n939_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n905_), .ZN(new_n950_));
  AOI21_X1  g749(.A(KEYINPUT115), .B1(new_n581_), .B2(new_n808_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n755_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT54), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n906_), .A2(new_n899_), .A3(new_n755_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n949_), .B1(new_n955_), .B2(new_n898_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n956_), .A2(new_n957_), .A3(new_n709_), .A4(new_n941_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n909_), .A2(new_n709_), .A3(new_n939_), .A4(new_n941_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(KEYINPUT119), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n958_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(new_n958_), .B2(new_n960_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n962_), .A2(new_n963_), .A3(new_n315_), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n959_), .A2(KEYINPUT119), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n959_), .A2(KEYINPUT119), .ZN(new_n966_));
  OAI21_X1  g765(.A(KEYINPUT61), .B1(new_n965_), .B2(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n958_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n968_));
  AOI21_X1  g767(.A(G155gat), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n964_), .A2(new_n969_), .ZN(G1346gat));
  NAND3_X1  g769(.A1(new_n943_), .A2(new_n316_), .A3(new_n707_), .ZN(new_n971_));
  NOR3_X1   g770(.A1(new_n940_), .A2(new_n755_), .A3(new_n942_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n316_), .B2(new_n972_), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT120), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n973_), .B(new_n974_), .ZN(G1347gat));
  AOI21_X1  g774(.A(new_n352_), .B1(new_n955_), .B2(new_n898_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n782_), .A2(new_n484_), .A3(new_n378_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n220_), .B1(new_n979_), .B2(new_n710_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n981_));
  OR2_X1    g780(.A1(new_n980_), .A2(new_n981_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n979_), .A2(new_n710_), .A3(new_n213_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n980_), .A2(new_n981_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n982_), .A2(new_n983_), .A3(new_n984_), .ZN(G1348gat));
  NAND2_X1  g784(.A1(new_n979_), .A2(new_n586_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n986_), .A2(new_n216_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n987_), .B1(new_n212_), .B2(new_n986_), .ZN(G1349gat));
  NOR2_X1   g787(.A1(new_n978_), .A2(new_n700_), .ZN(new_n989_));
  MUX2_X1   g788(.A(G183gat), .B(new_n238_), .S(new_n989_), .Z(G1350gat));
  NAND3_X1  g789(.A1(new_n707_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n991_));
  XOR2_X1   g790(.A(new_n991_), .B(KEYINPUT122), .Z(new_n992_));
  NAND2_X1  g791(.A1(new_n979_), .A2(new_n992_), .ZN(new_n993_));
  OAI21_X1  g792(.A(G190gat), .B1(new_n978_), .B2(new_n755_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n993_), .A2(new_n994_), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n995_), .B(KEYINPUT123), .ZN(G1351gat));
  NOR3_X1   g795(.A1(new_n940_), .A2(new_n378_), .A3(new_n782_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n997_), .A2(new_n710_), .ZN(new_n998_));
  AND3_X1   g797(.A1(new_n998_), .A2(KEYINPUT124), .A3(new_n278_), .ZN(new_n999_));
  AOI21_X1  g798(.A(KEYINPUT124), .B1(new_n998_), .B2(new_n278_), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(new_n998_), .A2(new_n278_), .ZN(new_n1001_));
  NOR3_X1   g800(.A1(new_n999_), .A2(new_n1000_), .A3(new_n1001_), .ZN(G1352gat));
  OAI21_X1  g801(.A(KEYINPUT126), .B1(new_n281_), .B2(KEYINPUT125), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1003_), .B1(KEYINPUT126), .B2(new_n281_), .ZN(new_n1004_));
  NAND3_X1  g803(.A1(new_n956_), .A2(new_n379_), .A3(new_n783_), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n1005_), .A2(new_n924_), .ZN(new_n1006_));
  MUX2_X1   g805(.A(new_n1003_), .B(new_n1004_), .S(new_n1006_), .Z(G1353gat));
  NAND2_X1  g806(.A1(new_n997_), .A2(new_n709_), .ZN(new_n1008_));
  NOR2_X1   g807(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1009_));
  AND2_X1   g808(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1010_));
  NOR3_X1   g809(.A1(new_n1008_), .A2(new_n1009_), .A3(new_n1010_), .ZN(new_n1011_));
  AOI21_X1  g810(.A(new_n1011_), .B1(new_n1008_), .B2(new_n1009_), .ZN(G1354gat));
  NAND3_X1  g811(.A1(new_n997_), .A2(new_n285_), .A3(new_n707_), .ZN(new_n1013_));
  OAI21_X1  g812(.A(G218gat), .B1(new_n1005_), .B2(new_n755_), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n1013_), .A2(new_n1014_), .ZN(G1355gat));
endmodule


