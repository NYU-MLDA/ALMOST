//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_;
  XNOR2_X1  g000(.A(KEYINPUT5), .B(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G204gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G120gat), .B(G148gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT66), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n208_), .A2(KEYINPUT9), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(KEYINPUT9), .B2(new_n208_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT10), .B(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(new_n214_), .A3(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n214_), .B1(new_n213_), .B2(G106gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n212_), .A2(new_n215_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n209_), .A2(new_n210_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n207_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT68), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n227_), .A3(new_n207_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n231_), .A2(new_n217_), .A3(new_n218_), .A4(KEYINPUT67), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n233_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n232_), .A2(new_n219_), .A3(new_n234_), .A4(new_n220_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n229_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n230_), .B1(new_n229_), .B2(new_n235_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n223_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n223_), .B(KEYINPUT69), .C1(new_n236_), .C2(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G78gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n244_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n246_), .B1(new_n249_), .B2(new_n245_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n240_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT64), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n238_), .A2(KEYINPUT12), .A3(new_n250_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n259_), .A2(new_n252_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n206_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n257_), .A2(new_n262_), .A3(new_n206_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(KEYINPUT70), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT70), .B1(new_n264_), .B2(new_n265_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT13), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT13), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G64gat), .B(G92gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G197gat), .B(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n283_));
  OR2_X1    g082(.A1(G211gat), .A2(G218gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G211gat), .A2(G218gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G197gat), .B(G204gat), .Z(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(KEYINPUT21), .B2(new_n282_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT24), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT78), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n297_));
  AND2_X1   g096(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n299_));
  OAI22_X1  g098(.A1(new_n296_), .A2(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G169gat), .ZN(new_n301_));
  INV_X1    g100(.A(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(KEYINPUT24), .A4(new_n292_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n295_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT79), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT23), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n303_), .A2(KEYINPUT24), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT79), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n295_), .A2(new_n300_), .A3(new_n312_), .A4(new_n305_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT80), .B(G176gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT22), .B(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n308_), .B(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n317_), .B(new_n292_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n291_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n303_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n309_), .A2(new_n310_), .A3(new_n300_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n288_), .A2(new_n290_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n326_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n322_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n314_), .A2(new_n321_), .A3(new_n291_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n323_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n326_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n280_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G127gat), .A2(G134gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G127gat), .ZN(new_n344_));
  INV_X1    g143(.A(G134gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT82), .B1(new_n346_), .B2(new_n339_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n338_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n342_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(KEYINPUT82), .A3(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n337_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT85), .B1(new_n358_), .B2(KEYINPUT1), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  AND2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n357_), .B1(new_n362_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  INV_X1    g167(.A(G141gat), .ZN(new_n369_));
  INV_X1    g168(.A(G148gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n353_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .A4(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n363_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n358_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n352_), .B1(new_n367_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n366_), .A2(new_n381_), .A3(new_n359_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n356_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n376_), .A2(new_n377_), .A3(new_n358_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n383_), .A2(new_n351_), .A3(new_n348_), .A4(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n379_), .A2(KEYINPUT4), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n384_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n352_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(new_n209_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT0), .B(G57gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n393_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n391_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n402_), .B2(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n314_), .A2(new_n321_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n323_), .B1(new_n405_), .B2(new_n330_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n329_), .A2(KEYINPUT90), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n329_), .A2(KEYINPUT90), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n291_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n326_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n333_), .A2(new_n334_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(new_n325_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n280_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n336_), .A2(new_n404_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n278_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n325_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n405_), .A2(new_n330_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n331_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT20), .A3(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n419_), .A3(new_n279_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n415_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n386_), .A2(new_n391_), .A3(new_n389_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n379_), .A2(new_n392_), .A3(new_n385_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n398_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n403_), .A2(KEYINPUT33), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n430_), .B(new_n397_), .C1(new_n402_), .C2(new_n399_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n414_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n387_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G22gat), .B(G50gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT28), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n436_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n330_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT86), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT87), .B(KEYINPUT29), .Z(new_n446_));
  OAI211_X1 g245(.A(new_n330_), .B(new_n445_), .C1(new_n434_), .C2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G78gat), .B(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n440_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n444_), .A2(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n448_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n439_), .A3(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT91), .B1(new_n433_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n279_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n332_), .A2(new_n335_), .A3(new_n278_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT89), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n429_), .A2(new_n431_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n415_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n427_), .A4(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n336_), .A2(new_n404_), .A3(new_n413_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n452_), .A2(new_n456_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n415_), .A2(new_n420_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n420_), .A2(KEYINPUT93), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n278_), .B(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n416_), .A2(new_n419_), .A3(new_n477_), .A4(new_n279_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n472_), .B1(new_n479_), .B2(KEYINPUT27), .ZN(new_n480_));
  INV_X1    g279(.A(new_n404_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT94), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(KEYINPUT27), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n471_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n486_));
  INV_X1    g285(.A(new_n482_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n458_), .A2(new_n469_), .A3(new_n483_), .A4(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G15gat), .B(G43gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT30), .B(G99gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(G71gat), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n314_), .A2(new_n321_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n492_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n348_), .A2(KEYINPUT31), .A3(new_n351_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT31), .B1(new_n348_), .B2(new_n351_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT81), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n405_), .A2(new_n494_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n502_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n490_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT83), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n502_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n497_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n491_), .B1(new_n503_), .B2(new_n496_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n490_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n505_), .A3(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n508_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT83), .B1(new_n508_), .B2(new_n516_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT84), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n516_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n514_), .B2(new_n505_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n509_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n404_), .B1(new_n519_), .B2(new_n525_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n480_), .A2(new_n457_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n489_), .A2(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT71), .B(G15gat), .ZN(new_n531_));
  INV_X1    g330(.A(G22gat), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G1gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n532_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G1gat), .B(G8gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G29gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT15), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(KEYINPUT76), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(KEYINPUT76), .B2(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n540_), .B(new_n546_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT77), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n273_), .A2(new_n530_), .A3(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT74), .ZN(new_n567_));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(KEYINPUT72), .A3(KEYINPUT17), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n540_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n250_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n574_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT75), .Z(new_n582_));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n242_), .A2(new_n543_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT34), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n238_), .A2(new_n544_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n585_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  OAI211_X1 g394(.A(new_n584_), .B(new_n589_), .C1(new_n585_), .C2(new_n588_), .ZN(new_n596_));
  AND4_X1   g395(.A1(new_n583_), .A2(new_n592_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n595_), .B(KEYINPUT36), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n582_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n565_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT95), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n534_), .A3(new_n404_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n564_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n272_), .A2(new_n612_), .A3(new_n581_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n601_), .B1(new_n613_), .B2(KEYINPUT96), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n489_), .A2(new_n527_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT84), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n523_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n481_), .B(new_n529_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n614_), .B(new_n619_), .C1(KEYINPUT96), .C2(new_n613_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n481_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n609_), .A2(new_n610_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n621_), .A3(new_n622_), .ZN(G1324gat));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n620_), .A2(new_n485_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT39), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n608_), .A2(new_n535_), .A3(new_n480_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n625_), .B2(G8gat), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n628_), .B(new_n624_), .C1(new_n630_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n629_), .A2(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n620_), .B2(new_n527_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT98), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(G15gat), .C1(new_n620_), .C2(new_n527_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n608_), .A2(new_n643_), .A3(new_n526_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n637_), .A2(KEYINPUT41), .A3(new_n639_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n642_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT99), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n642_), .A2(new_n644_), .A3(new_n648_), .A4(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n620_), .B2(new_n468_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n468_), .A2(G22gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT100), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n608_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT91), .B(new_n457_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n486_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n480_), .A2(KEYINPUT94), .A3(new_n482_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n526_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n618_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n657_), .B(new_n605_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n605_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n530_), .B2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n619_), .A2(KEYINPUT101), .A3(new_n657_), .A4(new_n605_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n582_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n273_), .A2(new_n564_), .A3(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n672_), .A2(new_n677_), .A3(new_n674_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT104), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n672_), .A2(new_n677_), .A3(new_n674_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT104), .B(new_n682_), .C1(new_n684_), .C2(new_n678_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n404_), .B(new_n676_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n684_), .B2(new_n678_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n675_), .B1(new_n692_), .B2(new_n685_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(KEYINPUT105), .A3(new_n404_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(G29gat), .A3(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n673_), .A2(new_n602_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n565_), .A2(new_n696_), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n697_), .A2(G29gat), .A3(new_n481_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n693_), .B2(new_n480_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n485_), .A2(G36gat), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n697_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n697_), .B2(new_n705_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n700_), .B1(new_n702_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n708_), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n485_), .B(new_n675_), .C1(new_n692_), .C2(new_n685_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT46), .B(new_n710_), .C1(new_n711_), .C2(new_n701_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1329gat));
  NAND2_X1  g512(.A1(new_n526_), .A2(G43gat), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n675_), .B(new_n714_), .C1(new_n692_), .C2(new_n685_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT107), .B(G43gat), .Z(new_n718_));
  INV_X1    g517(.A(new_n697_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n526_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n717_), .A3(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT47), .B1(new_n715_), .B2(new_n720_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n719_), .B2(new_n457_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n457_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n693_), .B2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n272_), .A2(new_n612_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n619_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n606_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n404_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n602_), .A3(new_n673_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n481_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(G57gat), .B2(new_n735_), .ZN(G1332gat));
  OR3_X1    g535(.A1(new_n731_), .A2(G64gat), .A3(new_n485_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G64gat), .B1(new_n734_), .B2(new_n485_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT48), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT48), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(G1333gat));
  OR3_X1    g540(.A1(new_n731_), .A2(G71gat), .A3(new_n527_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n734_), .A2(new_n527_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(G71gat), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G71gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1334gat));
  OR3_X1    g546(.A1(new_n731_), .A2(G78gat), .A3(new_n468_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G78gat), .B1(new_n734_), .B2(new_n468_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT50), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT50), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(G1335gat));
  NAND2_X1  g551(.A1(new_n730_), .A2(new_n696_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n209_), .A3(new_n404_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n672_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n272_), .A2(new_n612_), .A3(new_n673_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT109), .B1(new_n756_), .B2(new_n758_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n481_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n755_), .B1(new_n763_), .B2(new_n209_), .ZN(G1336gat));
  AOI21_X1  g563(.A(G92gat), .B1(new_n754_), .B2(new_n480_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n762_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n485_), .A2(new_n210_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT110), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n765_), .B1(new_n766_), .B2(new_n768_), .ZN(G1337gat));
  NOR3_X1   g568(.A1(new_n753_), .A2(new_n213_), .A3(new_n527_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n759_), .A2(new_n526_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G99gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n772_), .B(new_n773_), .Z(G1338gat));
  NAND3_X1  g573(.A1(new_n672_), .A2(new_n457_), .A3(new_n757_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT113), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n672_), .A2(new_n777_), .A3(new_n757_), .A4(new_n457_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(G106gat), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n776_), .A2(KEYINPUT114), .A3(G106gat), .A4(new_n778_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(KEYINPUT52), .A3(new_n782_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n753_), .A2(G106gat), .A3(new_n468_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT112), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n779_), .A2(new_n780_), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n272_), .A2(new_n564_), .A3(new_n606_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n790_), .B(new_n791_), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n259_), .A2(new_n252_), .A3(new_n261_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT116), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n259_), .A2(new_n252_), .A3(new_n795_), .A4(new_n261_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n256_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n794_), .A2(new_n799_), .A3(new_n256_), .A4(new_n796_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n262_), .B(KEYINPUT55), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n205_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT119), .A3(new_n806_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(KEYINPUT119), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n551_), .A2(new_n554_), .A3(new_n562_), .ZN(new_n809_));
  MUX2_X1   g608(.A(new_n552_), .B(new_n549_), .S(new_n553_), .Z(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n562_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n265_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(new_n808_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n807_), .A2(new_n808_), .A3(KEYINPUT58), .A4(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n605_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n561_), .A2(new_n563_), .A3(new_n265_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n269_), .A2(new_n811_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT57), .B(new_n602_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT118), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n602_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(KEYINPUT118), .A3(new_n827_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n816_), .A2(KEYINPUT120), .A3(new_n605_), .A4(new_n817_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n820_), .A2(new_n829_), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n581_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n792_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n526_), .A2(new_n404_), .A3(new_n529_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n818_), .A2(new_n828_), .A3(new_n824_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n582_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n790_), .B(new_n791_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n839_), .A2(new_n840_), .B1(KEYINPUT121), .B2(new_n836_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n837_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n832_), .A2(new_n833_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n840_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n836_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(KEYINPUT59), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n839_), .A2(new_n840_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n842_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n835_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n844_), .A2(new_n854_), .A3(G113gat), .A4(new_n612_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n834_), .A2(new_n836_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n858_), .B2(new_n564_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n855_), .A2(new_n859_), .ZN(G1340gat));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT123), .B(G120gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n272_), .B2(KEYINPUT60), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n857_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n861_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n861_), .A2(new_n857_), .A3(new_n867_), .A4(new_n864_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n272_), .B1(new_n848_), .B2(new_n852_), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n868_), .A2(new_n869_), .B1(new_n863_), .B2(new_n870_), .ZN(G1341gat));
  XOR2_X1   g670(.A(KEYINPUT125), .B(G127gat), .Z(new_n872_));
  NAND4_X1  g671(.A1(new_n844_), .A2(new_n854_), .A3(new_n581_), .A4(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n344_), .B1(new_n858_), .B2(new_n582_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  NAND4_X1  g674(.A1(new_n844_), .A2(new_n854_), .A3(G134gat), .A4(new_n605_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n345_), .B1(new_n858_), .B2(new_n602_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n834_), .A2(new_n481_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n480_), .A2(new_n468_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n612_), .A3(new_n527_), .A4(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g681(.A1(new_n879_), .A2(new_n273_), .A3(new_n527_), .A4(new_n880_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g683(.A1(new_n879_), .A2(new_n527_), .A3(new_n673_), .A4(new_n880_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  AND4_X1   g686(.A1(G162gat), .A2(new_n879_), .A3(new_n527_), .A4(new_n880_), .ZN(new_n888_));
  INV_X1    g687(.A(G162gat), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n879_), .A2(new_n527_), .A3(new_n601_), .A4(new_n880_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n605_), .B1(new_n889_), .B2(new_n890_), .ZN(G1347gat));
  NAND2_X1  g690(.A1(new_n528_), .A2(new_n480_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n457_), .B(new_n892_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n301_), .B1(new_n893_), .B2(new_n612_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT62), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n893_), .B(KEYINPUT126), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n612_), .A3(new_n316_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1348gat));
  NAND2_X1  g697(.A1(new_n846_), .A2(new_n468_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n899_), .A2(new_n302_), .A3(new_n272_), .A4(new_n892_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n273_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n315_), .ZN(G1349gat));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n893_), .B(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n833_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n297_), .A2(new_n296_), .ZN(new_n906_));
  INV_X1    g705(.A(G183gat), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n899_), .A2(new_n582_), .A3(new_n892_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n905_), .A2(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n904_), .B2(new_n669_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n601_), .B1(new_n299_), .B2(new_n298_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n904_), .B2(new_n911_), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n834_), .A2(new_n485_), .A3(new_n526_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n612_), .A3(new_n487_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n273_), .A3(new_n487_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g716(.A1(new_n913_), .A2(new_n487_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT63), .B(G211gat), .Z(new_n919_));
  NAND3_X1  g718(.A1(new_n918_), .A2(new_n581_), .A3(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n913_), .A2(new_n487_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n833_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n920_), .A2(new_n923_), .ZN(G1354gat));
  AOI21_X1  g723(.A(new_n526_), .B1(new_n845_), .B2(new_n840_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n925_), .A2(new_n480_), .A3(new_n487_), .A4(new_n601_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT127), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n913_), .A2(new_n928_), .A3(new_n487_), .A4(new_n601_), .ZN(new_n929_));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n918_), .A2(G218gat), .A3(new_n605_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1355gat));
endmodule


