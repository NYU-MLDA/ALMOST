//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n975_, new_n976_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n986_, new_n987_, new_n988_, new_n990_, new_n991_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G1gat), .A2(G8gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT14), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G1gat), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(new_n203_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n202_), .A2(new_n203_), .A3(new_n208_), .A4(new_n204_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G231gat), .A2(G233gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n212_), .B(new_n213_), .Z(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT71), .B(G71gat), .ZN(new_n215_));
  INV_X1    g014(.A(G78gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G57gat), .B(G64gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n215_), .A2(new_n216_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n216_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n219_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n221_), .B(new_n222_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n214_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G155gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT16), .ZN(new_n230_));
  XOR2_X1   g029(.A(G183gat), .B(G211gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(KEYINPUT17), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n227_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT76), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G232gat), .A2(G233gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT34), .Z(new_n238_));
  INV_X1    g037(.A(KEYINPUT35), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT73), .Z(new_n241_));
  NAND2_X1  g040(.A1(G99gat), .A2(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT6), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G99gat), .A3(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n245_), .A3(KEYINPUT68), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT67), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n258_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n261_));
  NOR2_X1   g060(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n262_));
  INV_X1    g061(.A(G85gat), .ZN(new_n263_));
  INV_X1    g062(.A(G92gat), .ZN(new_n264_));
  OAI22_X1  g063(.A1(new_n261_), .A2(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n264_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n260_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT69), .B1(new_n255_), .B2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n243_), .A2(new_n245_), .A3(KEYINPUT68), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT68), .B1(new_n243_), .B2(new_n245_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .A4(new_n253_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G85gat), .B(G92gat), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT8), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n248_), .A2(new_n254_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT7), .ZN(new_n280_));
  INV_X1    g079(.A(G99gat), .ZN(new_n281_));
  INV_X1    g080(.A(G106gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n278_), .B1(new_n279_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n285_), .A2(new_n287_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(KEYINPUT70), .A3(new_n284_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n277_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT8), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n286_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n275_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT15), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G43gat), .B(G50gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(new_n296_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n294_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G29gat), .B(G36gat), .Z(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n296_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT15), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n241_), .B1(new_n293_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n307_));
  INV_X1    g106(.A(new_n284_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n287_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n246_), .A3(new_n289_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n276_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT8), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n313_), .A2(new_n286_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n302_), .A2(new_n303_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n307_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND4_X1   g115(.A1(new_n307_), .A2(new_n275_), .A3(new_n292_), .A4(new_n315_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n306_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n238_), .A2(new_n239_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n321_), .B(new_n306_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G190gat), .B(G218gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G134gat), .B(G162gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT36), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT74), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n325_), .B(KEYINPUT36), .Z(new_n329_));
  INV_X1    g128(.A(new_n315_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n293_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n314_), .A2(new_n307_), .A3(new_n315_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n321_), .B1(new_n333_), .B2(new_n306_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n322_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n329_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n320_), .A2(new_n337_), .A3(new_n322_), .A4(new_n326_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n328_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT37), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT37), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n327_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n320_), .A2(new_n322_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(KEYINPUT75), .A3(new_n329_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n236_), .B1(new_n340_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT77), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n351_));
  INV_X1    g150(.A(G141gat), .ZN(new_n352_));
  INV_X1    g151(.A(G148gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT3), .ZN(new_n355_));
  NOR3_X1   g154(.A1(KEYINPUT88), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n355_), .A2(new_n358_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G155gat), .B(G162gat), .Z(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n359_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n363_), .A2(new_n364_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n373_), .A2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT94), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n373_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n375_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n372_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n375_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n364_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n361_), .A2(new_n362_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n357_), .B1(new_n367_), .B2(new_n351_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n389_), .B2(new_n358_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n370_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT94), .B(new_n385_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n384_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n384_), .B2(new_n392_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n394_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n376_), .A2(new_n377_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n401_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n403_), .B1(new_n405_), .B2(new_n372_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n395_), .B(new_n400_), .C1(new_n402_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n393_), .A2(KEYINPUT4), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n408_), .A2(new_n409_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n410_), .B2(new_n400_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  NOR3_X1   g211(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(KEYINPUT93), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n417_));
  INV_X1    g216(.A(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n413_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n423_));
  INV_X1    g222(.A(G183gat), .ZN(new_n424_));
  INV_X1    g223(.A(G190gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n416_), .A2(new_n419_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT24), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n422_), .A2(new_n423_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT24), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT92), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n439_), .A3(KEYINPUT24), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441_));
  INV_X1    g240(.A(G169gat), .ZN(new_n442_));
  INV_X1    g241(.A(G176gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n444_), .A3(new_n430_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n433_), .B(new_n434_), .C1(new_n438_), .C2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n425_), .A2(KEYINPUT26), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT26), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G190gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n424_), .A2(KEYINPUT25), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT25), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(G183gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT91), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(G183gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n424_), .A2(KEYINPUT25), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n450_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n428_), .B1(new_n446_), .B2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G197gat), .A2(G204gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G197gat), .A2(G204gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT21), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT21), .ZN(new_n465_));
  INV_X1    g264(.A(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(new_n461_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G211gat), .B(G218gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G211gat), .B(G218gat), .Z(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(KEYINPUT21), .A3(new_n462_), .A4(new_n463_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n412_), .B1(new_n460_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n469_), .A2(new_n471_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT25), .B1(new_n424_), .B2(KEYINPUT81), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n452_), .A3(G183gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n478_), .A2(new_n480_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n429_), .B1(G169gat), .B2(G176gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(new_n444_), .A3(new_n430_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n433_), .A2(new_n481_), .A3(new_n483_), .A4(new_n434_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n427_), .A2(KEYINPUT83), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n422_), .A2(new_n426_), .A3(new_n486_), .A4(new_n423_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n418_), .A2(new_n413_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n477_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n473_), .A2(new_n476_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n450_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n458_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n457_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n437_), .A2(new_n444_), .A3(new_n430_), .A4(new_n440_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n422_), .A2(new_n423_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n444_), .A2(new_n430_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(new_n429_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n477_), .A3(new_n428_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n484_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n472_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT20), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n491_), .B1(new_n504_), .B2(new_n476_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G8gat), .B(G36gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT18), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT32), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n505_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n460_), .A2(new_n472_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(KEYINPUT20), .A3(new_n490_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n475_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT20), .A4(new_n476_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n411_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT96), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT33), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n407_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n408_), .A2(new_n409_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n400_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n522_), .A2(new_n524_), .A3(KEYINPUT96), .A4(KEYINPUT33), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n395_), .A2(new_n400_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n402_), .A2(new_n406_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n515_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n509_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n516_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n476_), .B1(new_n473_), .B2(new_n490_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n400_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n394_), .B1(new_n405_), .B2(new_n372_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n402_), .B2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n530_), .A2(new_n531_), .A3(new_n535_), .A4(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n518_), .B1(new_n526_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G78gat), .B(G106gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n372_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT28), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n543_), .A2(KEYINPUT28), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n541_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n543_), .A2(KEYINPUT28), .ZN(new_n548_));
  INV_X1    g347(.A(new_n541_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n472_), .B1(new_n372_), .B2(new_n542_), .ZN(new_n552_));
  AND2_X1   g351(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n553_));
  NOR2_X1   g352(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(G228gat), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(KEYINPUT90), .A3(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(KEYINPUT90), .Z(new_n557_));
  OAI211_X1 g356(.A(new_n472_), .B(new_n557_), .C1(new_n372_), .C2(new_n542_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G22gat), .B(G50gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n551_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n565_), .A2(new_n550_), .A3(new_n547_), .A4(new_n561_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n540_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n411_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n505_), .A2(new_n532_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT27), .A3(new_n531_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT98), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n535_), .A2(new_n531_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT27), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AOI211_X1 g374(.A(KEYINPUT98), .B(KEYINPUT27), .C1(new_n535_), .C2(new_n531_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n569_), .B(new_n571_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n568_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G227gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(G71gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G15gat), .B(G43gat), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT85), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(G99gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n583_), .B(KEYINPUT85), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n281_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n582_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(G99gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n281_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n581_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n502_), .B(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n385_), .B(KEYINPUT31), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n595_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n601_), .A2(KEYINPUT86), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(KEYINPUT86), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n597_), .A2(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI221_X1 g405(.A(new_n600_), .B1(new_n598_), .B2(new_n597_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n567_), .B(new_n571_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n411_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n578_), .A2(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT64), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n275_), .A2(new_n292_), .A3(new_n226_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n226_), .B1(new_n275_), .B2(new_n292_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n615_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n226_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n293_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n275_), .A2(new_n292_), .A3(new_n226_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n615_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT5), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n622_), .A2(new_n627_), .A3(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n624_), .A2(KEYINPUT12), .A3(new_n625_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n614_), .B1(new_n634_), .B2(new_n620_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n635_), .B2(new_n626_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(new_n636_), .A3(KEYINPUT13), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT13), .B1(new_n633_), .B2(new_n636_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G169gat), .B(G197gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(new_n642_), .Z(new_n643_));
  INV_X1    g442(.A(new_n211_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n202_), .A2(new_n204_), .B1(new_n203_), .B2(new_n208_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n303_), .B(new_n302_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n315_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n299_), .A2(new_n212_), .A3(new_n304_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT78), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n649_), .A4(new_n647_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n649_), .A3(new_n647_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT78), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n643_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT79), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n657_), .A2(new_n651_), .A3(new_n654_), .A4(new_n643_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT80), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT80), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n655_), .A2(new_n663_), .A3(new_n657_), .A4(new_n643_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n660_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n640_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n612_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n350_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n206_), .A3(new_n411_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT38), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n640_), .A2(KEYINPUT99), .A3(new_n666_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n345_), .A2(new_n347_), .A3(new_n327_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n612_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n236_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n675_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n411_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT100), .A3(G1gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT100), .B1(new_n680_), .B2(G1gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n671_), .B1(new_n681_), .B2(new_n682_), .ZN(G1324gat));
  INV_X1    g482(.A(new_n571_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n533_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n509_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n574_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT98), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n573_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n684_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n669_), .A2(new_n207_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT39), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n679_), .A2(new_n691_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G8gat), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT39), .B(new_n207_), .C1(new_n679_), .C2(new_n691_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n697_), .B(new_n698_), .Z(G1325gat));
  INV_X1    g498(.A(G15gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n608_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n669_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n679_), .A2(new_n701_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n703_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(new_n703_), .B2(G15gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT102), .Z(G1326gat));
  INV_X1    g506(.A(G22gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n567_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n669_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n679_), .A2(new_n709_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G22gat), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(KEYINPUT42), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(KEYINPUT42), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1327gat));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n340_), .A2(new_n717_), .A3(new_n348_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT105), .B1(new_n612_), .B2(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n340_), .A2(new_n717_), .A3(new_n348_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n611_), .A2(new_n567_), .A3(new_n690_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n690_), .A2(new_n569_), .B1(new_n540_), .B2(new_n567_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n701_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n327_), .A2(KEYINPUT74), .B1(new_n346_), .B2(new_n329_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n341_), .B1(new_n727_), .B2(new_n338_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT75), .B1(new_n346_), .B2(new_n329_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n329_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n344_), .B(new_n730_), .C1(new_n320_), .C2(new_n322_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n729_), .A2(new_n731_), .A3(new_n342_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n726_), .B1(new_n728_), .B2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n340_), .A2(KEYINPUT104), .A3(new_n348_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n719_), .A2(new_n725_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n675_), .A2(new_n236_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n716_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n725_), .A2(new_n719_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(new_n736_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n738_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(KEYINPUT44), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n411_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G29gat), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n676_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n678_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n668_), .A2(new_n749_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n746_), .A2(G29gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1328gat));
  OR2_X1    g551(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n750_), .A2(G36gat), .A3(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT45), .Z(new_n757_));
  NAND3_X1  g556(.A1(new_n739_), .A2(new_n744_), .A3(new_n691_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(KEYINPUT106), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n739_), .A2(new_n744_), .A3(new_n760_), .A4(new_n691_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G36gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT46), .B(new_n757_), .C1(new_n759_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1329gat));
  NAND4_X1  g566(.A1(new_n739_), .A2(new_n744_), .A3(G43gat), .A4(new_n701_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n750_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G43gat), .B1(new_n769_), .B2(new_n701_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(KEYINPUT108), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(KEYINPUT108), .B2(new_n768_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n773_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n771_), .B(new_n775_), .C1(KEYINPUT108), .C2(new_n768_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1330gat));
  INV_X1    g576(.A(G50gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n750_), .B2(new_n567_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n567_), .A2(new_n778_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n745_), .B2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT110), .Z(G1331gat));
  NOR3_X1   g582(.A1(new_n612_), .A2(new_n666_), .A3(new_n640_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n350_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(G57gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n411_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n640_), .A2(new_n666_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n677_), .A2(new_n678_), .A3(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT111), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(new_n411_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n792_), .B2(new_n787_), .ZN(G1332gat));
  INV_X1    g592(.A(G64gat), .ZN(new_n794_));
  INV_X1    g593(.A(new_n755_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT48), .Z(new_n797_));
  NAND3_X1  g596(.A1(new_n786_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1333gat));
  NAND3_X1  g598(.A1(new_n786_), .A2(new_n580_), .A3(new_n701_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n580_), .B1(new_n791_), .B2(new_n701_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(G1334gat));
  AOI21_X1  g604(.A(new_n216_), .B1(new_n791_), .B2(new_n709_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT50), .Z(new_n807_));
  NAND3_X1  g606(.A1(new_n786_), .A2(new_n216_), .A3(new_n709_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1335gat));
  NAND2_X1  g608(.A1(new_n784_), .A2(new_n749_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n263_), .A3(new_n411_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n742_), .A2(new_n236_), .A3(new_n789_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(new_n411_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(new_n263_), .ZN(G1336gat));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n264_), .A3(new_n691_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n813_), .A2(new_n795_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n264_), .ZN(G1337gat));
  AND4_X1   g617(.A1(new_n701_), .A2(new_n811_), .A3(new_n249_), .A4(new_n251_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n813_), .A2(new_n701_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G99gat), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g621(.A1(new_n811_), .A2(new_n709_), .A3(new_n250_), .A4(new_n252_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n742_), .A2(new_n709_), .A3(new_n236_), .A4(new_n789_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  AND4_X1   g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .A4(G106gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n282_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n825_), .A2(new_n828_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n823_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n823_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n609_), .A2(new_n746_), .A3(new_n608_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n633_), .A2(new_n636_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n643_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT115), .B1(new_n652_), .B2(new_n647_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n839_), .A2(new_n649_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n652_), .A2(KEYINPUT115), .A3(new_n647_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n665_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n837_), .A2(KEYINPUT116), .A3(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n666_), .A2(new_n633_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n634_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n622_), .A2(KEYINPUT55), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n632_), .B1(new_n635_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n854_), .A3(KEYINPUT56), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n850_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n748_), .B1(new_n849_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n844_), .A2(new_n633_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n852_), .A2(new_n854_), .A3(KEYINPUT56), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n855_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n729_), .A2(new_n731_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n867_), .A2(new_n343_), .B1(new_n339_), .B2(KEYINPUT37), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT58), .B(new_n862_), .C1(new_n863_), .C2(new_n855_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT116), .B1(new_n837_), .B2(new_n844_), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n846_), .B(new_n843_), .C1(new_n633_), .C2(new_n636_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n666_), .B(new_n633_), .C1(new_n863_), .C2(new_n855_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n676_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n870_), .B1(new_n875_), .B2(KEYINPUT57), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n861_), .B1(new_n876_), .B2(KEYINPUT117), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n870_), .B(new_n878_), .C1(new_n875_), .C2(KEYINPUT57), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n678_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT13), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n837_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n637_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n666_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n349_), .A2(new_n881_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT114), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n349_), .A2(new_n885_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT54), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n349_), .A2(new_n890_), .A3(new_n885_), .A4(new_n881_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n835_), .B(new_n836_), .C1(new_n880_), .C2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n836_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n236_), .B1(new_n876_), .B2(new_n861_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n892_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n894_), .B1(new_n835_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n666_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G113gat), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n892_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n836_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n899_), .A2(G113gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n902_), .B2(new_n903_), .ZN(G1340gat));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905_));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n640_), .B1(new_n902_), .B2(KEYINPUT59), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n894_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n640_), .B2(KEYINPUT60), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(KEYINPUT60), .B2(new_n906_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n902_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n905_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n836_), .A2(new_n835_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n877_), .A2(new_n879_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n236_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n915_), .B2(new_n892_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n884_), .B1(new_n897_), .B2(new_n835_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G120gat), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n911_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n918_), .A2(KEYINPUT118), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n912_), .A2(new_n920_), .ZN(G1341gat));
  OAI21_X1  g720(.A(G127gat), .B1(new_n898_), .B2(new_n236_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n236_), .A2(G127gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n902_), .B2(new_n923_), .ZN(G1342gat));
  NAND2_X1  g723(.A1(new_n340_), .A2(new_n348_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G134gat), .B1(new_n898_), .B2(new_n925_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n748_), .A2(G134gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n902_), .B2(new_n927_), .ZN(G1343gat));
  INV_X1    g727(.A(new_n901_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n755_), .A2(new_n411_), .A3(new_n709_), .A4(new_n608_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT119), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n666_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT120), .B(G141gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1344gat));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n884_), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT121), .B(G148gat), .Z(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1345gat));
  NAND2_X1  g737(.A1(new_n932_), .A2(new_n678_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1346gat));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n733_), .A2(new_n734_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n932_), .A2(G162gat), .A3(new_n943_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n929_), .A2(new_n748_), .A3(new_n931_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(G162gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n942_), .B1(new_n944_), .B2(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n932_), .A2(G162gat), .A3(new_n943_), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n948_), .B(KEYINPUT122), .C1(G162gat), .C2(new_n945_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1347gat));
  XOR2_X1   g749(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n795_), .A2(new_n611_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n709_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n666_), .B(new_n954_), .C1(new_n880_), .C2(new_n893_), .ZN(new_n955_));
  OAI211_X1 g754(.A(new_n442_), .B(new_n952_), .C1(new_n955_), .C2(KEYINPUT22), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n952_), .B1(new_n955_), .B2(KEYINPUT22), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n955_), .A2(new_n952_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n442_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n957_), .B1(new_n958_), .B2(new_n960_), .ZN(G1348gat));
  INV_X1    g760(.A(new_n954_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n915_), .B2(new_n892_), .ZN(new_n963_));
  AOI21_X1  g762(.A(G176gat), .B1(new_n963_), .B2(new_n884_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n901_), .A2(new_n567_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n953_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n966_), .A2(G176gat), .A3(new_n884_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n965_), .A2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(KEYINPUT124), .B1(new_n964_), .B2(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n954_), .B1(new_n880_), .B2(new_n893_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n443_), .B1(new_n970_), .B2(new_n640_), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n971_), .B(new_n972_), .C1(new_n965_), .C2(new_n967_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n969_), .A2(new_n973_), .ZN(G1349gat));
  NOR3_X1   g773(.A1(new_n236_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n975_));
  NAND4_X1  g774(.A1(new_n901_), .A2(new_n567_), .A3(new_n678_), .A4(new_n966_), .ZN(new_n976_));
  AOI22_X1  g775(.A1(new_n963_), .A2(new_n975_), .B1(new_n424_), .B2(new_n976_), .ZN(G1350gat));
  AOI21_X1  g776(.A(new_n425_), .B1(new_n963_), .B2(new_n868_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n676_), .A2(new_n492_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n970_), .A2(new_n979_), .ZN(new_n980_));
  OAI21_X1  g779(.A(KEYINPUT125), .B1(new_n978_), .B2(new_n980_), .ZN(new_n981_));
  OAI21_X1  g780(.A(G190gat), .B1(new_n970_), .B2(new_n925_), .ZN(new_n982_));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n982_), .B(new_n983_), .C1(new_n970_), .C2(new_n979_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n981_), .A2(new_n984_), .ZN(G1351gat));
  NAND3_X1  g784(.A1(new_n795_), .A2(new_n569_), .A3(new_n608_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n929_), .A2(new_n986_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n987_), .A2(new_n666_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g788(.A1(new_n987_), .A2(new_n884_), .ZN(new_n990_));
  INV_X1    g789(.A(G204gat), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n991_), .A2(KEYINPUT126), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n990_), .B(new_n992_), .ZN(G1353gat));
  NAND2_X1  g792(.A1(new_n987_), .A2(new_n678_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n995_));
  AND2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n994_), .A2(new_n995_), .A3(new_n996_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n997_), .B1(new_n994_), .B2(new_n995_), .ZN(G1354gat));
  INV_X1    g797(.A(G218gat), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n999_), .B1(new_n987_), .B2(new_n868_), .ZN(new_n1000_));
  INV_X1    g799(.A(new_n1000_), .ZN(new_n1001_));
  NOR4_X1   g800(.A1(new_n929_), .A2(G218gat), .A3(new_n748_), .A4(new_n986_), .ZN(new_n1002_));
  INV_X1    g801(.A(new_n1002_), .ZN(new_n1003_));
  NAND3_X1  g802(.A1(new_n1001_), .A2(KEYINPUT127), .A3(new_n1003_), .ZN(new_n1004_));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005_));
  OAI21_X1  g804(.A(new_n1005_), .B1(new_n1000_), .B2(new_n1002_), .ZN(new_n1006_));
  NAND2_X1  g805(.A1(new_n1004_), .A2(new_n1006_), .ZN(G1355gat));
endmodule


