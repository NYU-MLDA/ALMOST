//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT12), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212_));
  AND2_X1   g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n216_), .A2(new_n213_), .A3(new_n217_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n227_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(KEYINPUT64), .A3(new_n228_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n225_), .A2(new_n226_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n238_));
  NOR2_X1   g037(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n240_), .A2(new_n226_), .A3(new_n223_), .A4(new_n222_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n233_), .A2(new_n231_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n235_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n237_), .B(new_n215_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n242_), .B(new_n235_), .C1(new_n246_), .C2(new_n224_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT9), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n249_), .B2(new_n229_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n232_), .A2(KEYINPUT9), .A3(new_n228_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT10), .B(G99gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n251_), .C1(G106gat), .C2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n212_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n247_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n255_));
  AOI211_X1 g054(.A(KEYINPUT66), .B(new_n235_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n212_), .B(new_n253_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n211_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT12), .B1(new_n260_), .B2(new_n209_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n253_), .B(new_n208_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G230gat), .A2(G233gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n265_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n208_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(new_n263_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G176gat), .B(G204gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT69), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n266_), .A2(new_n278_), .A3(new_n269_), .A4(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n270_), .A2(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n284_), .A3(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G8gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT74), .B(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G43gat), .B(G50gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n290_), .A2(new_n295_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n287_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n299_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(KEYINPUT77), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n299_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n305_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G169gat), .B(G197gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT78), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G141gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n310_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n316_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n320_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n325_), .A3(KEYINPUT79), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n327_), .B(new_n320_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n286_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT92), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334_));
  INV_X1    g133(.A(G120gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT85), .B(G113gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(KEYINPUT2), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n347_), .B(new_n348_), .C1(new_n349_), .C2(new_n341_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n339_), .B(new_n340_), .C1(new_n344_), .C2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n343_), .A2(new_n345_), .ZN(new_n352_));
  AND3_X1   g151(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n339_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n333_), .B1(new_n338_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n338_), .A2(new_n357_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT4), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n332_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  INV_X1    g166(.A(G85gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT0), .B(G57gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n360_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT93), .B1(new_n373_), .B2(new_n332_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n366_), .B(new_n372_), .C1(new_n364_), .C2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n364_), .A2(new_n374_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n379_), .A2(KEYINPUT33), .A3(new_n372_), .A4(new_n366_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT84), .B(G176gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G169gat), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n381_), .A2(new_n382_), .B1(G169gat), .B2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(G183gat), .ZN(new_n384_));
  INV_X1    g183(.A(G190gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT23), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT83), .Z(new_n387_));
  OR3_X1    g186(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT23), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n383_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT24), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  MUX2_X1   g194(.A(new_n394_), .B(KEYINPUT24), .S(new_n395_), .Z(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n386_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT26), .B(G190gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT25), .B(G183gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n392_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G211gat), .B(G218gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(G197gat), .B(G204gat), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(KEYINPUT89), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n404_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(KEYINPUT21), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(KEYINPUT21), .B2(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(G183gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n397_), .B1(new_n411_), .B2(G190gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n383_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n398_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(KEYINPUT25), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT81), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(KEYINPUT82), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n384_), .B1(KEYINPUT82), .B2(new_n417_), .ZN(new_n419_));
  AOI211_X1 g218(.A(new_n414_), .B(new_n416_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n389_), .A2(new_n396_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n413_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n409_), .B(KEYINPUT20), .C1(new_n422_), .C2(new_n408_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n408_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n402_), .A2(new_n408_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT20), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432_));
  INV_X1    g231(.A(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT18), .B(G64gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n426_), .A2(new_n438_), .A3(new_n430_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n361_), .A2(new_n363_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n332_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n332_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n372_), .B1(new_n373_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT94), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(KEYINPUT94), .A3(new_n444_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n377_), .A2(new_n380_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n364_), .A2(new_n365_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n371_), .B1(new_n449_), .B2(new_n378_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n375_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n438_), .A2(KEYINPUT32), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n431_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT20), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n425_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(new_n425_), .B2(new_n423_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n351_), .A2(new_n356_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  XNOR2_X1  g262(.A(G22gat), .B(G50gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n461_), .B(new_n462_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n468_), .A3(KEYINPUT91), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G78gat), .B(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n465_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n408_), .B1(new_n459_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(G228gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(G228gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n408_), .B(new_n484_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n474_), .B(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n448_), .A2(new_n458_), .A3(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G71gat), .B(G99gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G43gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n422_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n338_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT30), .B(G15gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT31), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n494_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n492_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n456_), .A2(new_n436_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT27), .A3(new_n439_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT27), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n440_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n501_), .A2(new_n450_), .A3(new_n503_), .A4(new_n375_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n474_), .B(new_n486_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n499_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n489_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n503_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n451_), .A2(new_n498_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n331_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n300_), .B(new_n253_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n260_), .A2(KEYINPUT67), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n257_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n516_), .B2(new_n314_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT35), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G190gat), .B(G218gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n314_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n513_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n314_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n515_), .B2(new_n257_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n528_), .B(new_n532_), .C1(new_n535_), .C2(new_n514_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n522_), .B(new_n527_), .C1(new_n533_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT37), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n532_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT72), .B1(new_n517_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n536_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n544_), .B2(new_n522_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n522_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT73), .A3(new_n540_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n543_), .A2(new_n536_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n541_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n551_), .A3(new_n538_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n546_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n305_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n208_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT16), .B(G183gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n557_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n566_), .A2(KEYINPUT76), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(KEYINPUT76), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n554_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n512_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n291_), .A3(new_n451_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n569_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n552_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n512_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n451_), .ZN(new_n581_));
  OAI21_X1  g380(.A(G1gat), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n574_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n575_), .A2(new_n582_), .A3(new_n583_), .ZN(G1324gat));
  NAND3_X1  g383(.A1(new_n572_), .A2(new_n292_), .A3(new_n508_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n508_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G8gat), .B1(new_n580_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT95), .B(KEYINPUT40), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(G1325gat));
  OAI21_X1  g391(.A(G15gat), .B1(new_n580_), .B2(new_n498_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT41), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT41), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n571_), .A2(G15gat), .A3(new_n498_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(G1326gat));
  OR3_X1    g396(.A1(new_n571_), .A2(G22gat), .A3(new_n488_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G22gat), .B1(new_n580_), .B2(new_n488_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(KEYINPUT42), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(KEYINPUT42), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT96), .ZN(G1327gat));
  INV_X1    g402(.A(G29gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n576_), .A2(new_n330_), .A3(new_n286_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT43), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n507_), .A2(new_n511_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n554_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  AOI211_X1 g409(.A(KEYINPUT43), .B(new_n554_), .C1(new_n507_), .C2(new_n511_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT44), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT44), .B(new_n606_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n451_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n604_), .B1(new_n617_), .B2(KEYINPUT97), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(KEYINPUT97), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n569_), .A2(new_n552_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n512_), .A2(new_n604_), .A3(new_n451_), .A4(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(G1328gat));
  INV_X1    g421(.A(KEYINPUT46), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT98), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n508_), .A3(new_n615_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G36gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n512_), .A2(new_n620_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n627_), .A2(G36gat), .A3(new_n586_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT45), .Z(new_n629_));
  AOI21_X1  g428(.A(new_n624_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n623_), .A2(KEYINPUT98), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(G1329gat));
  NOR3_X1   g431(.A1(new_n627_), .A2(G43gat), .A3(new_n498_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n616_), .A2(new_n499_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n634_), .B2(G43gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g435(.A(G50gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n616_), .B2(new_n505_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n627_), .A2(G50gat), .A3(new_n488_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n638_), .A2(KEYINPUT99), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT99), .B1(new_n638_), .B2(new_n639_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1331gat));
  INV_X1    g441(.A(new_n286_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n329_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(new_n570_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G57gat), .B1(new_n646_), .B2(new_n451_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n578_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n451_), .A2(G57gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(G1332gat));
  INV_X1    g449(.A(G64gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n648_), .B2(new_n508_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT48), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n651_), .A3(new_n508_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1333gat));
  INV_X1    g454(.A(G71gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n646_), .A2(new_n656_), .A3(new_n499_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n648_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G71gat), .B1(new_n658_), .B2(new_n498_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT101), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(KEYINPUT101), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT100), .B(KEYINPUT49), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n663_), .B2(new_n664_), .ZN(G1334gat));
  INV_X1    g464(.A(G78gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n648_), .B2(new_n505_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT50), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n646_), .A2(new_n666_), .A3(new_n505_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1335gat));
  NOR2_X1   g469(.A1(new_n610_), .A2(new_n611_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n569_), .A3(new_n644_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n451_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n645_), .A2(new_n620_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n581_), .A2(G85gat), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n673_), .A2(G85gat), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT102), .Z(G1336gat));
  AOI21_X1  g476(.A(G92gat), .B1(new_n674_), .B2(new_n508_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n586_), .A2(new_n433_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n672_), .B2(new_n679_), .ZN(G1337gat));
  AOI21_X1  g479(.A(new_n220_), .B1(new_n672_), .B2(new_n499_), .ZN(new_n681_));
  AND2_X1   g480(.A1(KEYINPUT103), .A2(KEYINPUT51), .ZN(new_n682_));
  INV_X1    g481(.A(new_n252_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n674_), .A2(new_n683_), .A3(new_n499_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n681_), .A2(new_n682_), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(KEYINPUT103), .A2(KEYINPUT51), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT104), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n685_), .B(new_n687_), .ZN(G1338gat));
  NAND3_X1  g487(.A1(new_n674_), .A2(new_n221_), .A3(new_n505_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n644_), .A2(new_n569_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G106gat), .B1(new_n691_), .B2(new_n488_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT105), .B(KEYINPUT52), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n689_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT53), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n700_), .B(new_n689_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1339gat));
  OAI21_X1  g501(.A(new_n262_), .B1(new_n268_), .B2(KEYINPUT12), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n210_), .B1(new_n515_), .B2(new_n257_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(KEYINPUT55), .A4(new_n265_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n259_), .A2(new_n264_), .A3(KEYINPUT55), .A4(new_n265_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT107), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT55), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n259_), .A2(new_n264_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n267_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n266_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n707_), .B(new_n709_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(KEYINPUT56), .A4(new_n276_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n329_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n276_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT108), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n276_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n716_), .B(new_n717_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n309_), .A2(new_n310_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n315_), .A2(new_n311_), .A3(new_n307_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n320_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n322_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n322_), .B2(new_n724_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n577_), .B1(new_n721_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT57), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT57), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n714_), .A2(new_n276_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT56), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(KEYINPUT108), .A3(new_n718_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n716_), .A2(new_n717_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n729_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT110), .B(new_n734_), .C1(new_n740_), .C2(new_n577_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n728_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n714_), .A2(new_n743_), .A3(KEYINPUT56), .A4(new_n276_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n718_), .A2(KEYINPUT111), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n742_), .B(new_n744_), .C1(new_n745_), .C2(new_n720_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT58), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n554_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n737_), .A2(KEYINPUT111), .A3(new_n718_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n749_), .A2(KEYINPUT58), .A3(new_n744_), .A4(new_n742_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n733_), .A2(new_n741_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n576_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n330_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n570_), .B2(new_n755_), .ZN(new_n756_));
  AND4_X1   g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n554_), .A4(new_n569_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n753_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n509_), .A2(new_n499_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n451_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n581_), .B1(new_n753_), .B2(new_n759_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT112), .A3(new_n762_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n329_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT113), .B1(new_n768_), .B2(G113gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT112), .B1(new_n766_), .B2(new_n762_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n758_), .B1(new_n576_), .B2(new_n752_), .ZN(new_n771_));
  NOR4_X1   g570(.A1(new_n771_), .A2(new_n764_), .A3(new_n581_), .A4(new_n761_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n330_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  INV_X1    g573(.A(G113gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n763_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n771_), .A2(new_n581_), .A3(new_n761_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT59), .B1(new_n780_), .B2(KEYINPUT114), .ZN(new_n781_));
  OAI211_X1 g580(.A(G113gat), .B(new_n330_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n769_), .A2(new_n776_), .A3(new_n782_), .ZN(G1340gat));
  NAND2_X1  g582(.A1(new_n765_), .A2(new_n767_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n335_), .A2(KEYINPUT60), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n335_), .B1(new_n286_), .B2(KEYINPUT60), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n784_), .B(new_n788_), .C1(new_n787_), .C2(new_n786_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n779_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n781_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n286_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n789_), .B1(new_n792_), .B2(new_n335_), .ZN(G1341gat));
  AOI21_X1  g592(.A(G127gat), .B1(new_n784_), .B2(new_n569_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n791_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n569_), .A2(G127gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(G1342gat));
  AOI21_X1  g596(.A(G134gat), .B1(new_n784_), .B2(new_n577_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n609_), .A2(G134gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n795_), .B2(new_n799_), .ZN(G1343gat));
  NOR2_X1   g599(.A1(new_n488_), .A2(new_n499_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n508_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT110), .B1(new_n740_), .B2(new_n577_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n804_), .A2(KEYINPUT57), .B1(new_n750_), .B2(new_n748_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n569_), .B1(new_n805_), .B2(new_n741_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n451_), .B(new_n803_), .C1(new_n806_), .C2(new_n758_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n766_), .A2(KEYINPUT116), .A3(new_n803_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n330_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT117), .B(G141gat), .Z(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1344gat));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n643_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g615(.A(KEYINPUT61), .B(G155gat), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n811_), .B2(new_n569_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT118), .B(new_n576_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n818_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n766_), .B2(new_n803_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n803_), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n771_), .A2(new_n808_), .A3(new_n581_), .A4(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n569_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT118), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n811_), .A2(new_n819_), .A3(new_n569_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n817_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n822_), .A2(new_n829_), .ZN(G1346gat));
  NOR2_X1   g629(.A1(new_n552_), .A2(G162gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n554_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n833_));
  INV_X1    g632(.A(G162gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n832_), .B(new_n837_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1347gat));
  NAND2_X1  g638(.A1(new_n510_), .A2(new_n508_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n329_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT120), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n760_), .A2(new_n488_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G169gat), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(KEYINPUT62), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(KEYINPUT62), .ZN(new_n846_));
  INV_X1    g645(.A(new_n840_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n488_), .B(new_n847_), .C1(new_n806_), .C2(new_n758_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n760_), .A2(KEYINPUT121), .A3(new_n488_), .A4(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n330_), .A2(new_n382_), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n845_), .A2(new_n846_), .B1(new_n852_), .B2(new_n853_), .ZN(G1348gat));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n643_), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n381_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n848_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(G176gat), .A3(new_n643_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(KEYINPUT122), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1349gat));
  NOR3_X1   g662(.A1(new_n852_), .A2(new_n399_), .A3(new_n576_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n411_), .B1(new_n857_), .B2(new_n569_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1350gat));
  NAND3_X1  g665(.A1(new_n850_), .A2(new_n609_), .A3(new_n851_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n867_), .A2(new_n868_), .A3(G190gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n867_), .B2(G190gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n577_), .A2(new_n398_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT124), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n869_), .A2(new_n870_), .B1(new_n852_), .B2(new_n872_), .ZN(G1351gat));
  NOR3_X1   g672(.A1(new_n802_), .A2(new_n451_), .A3(new_n586_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n760_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n760_), .A2(KEYINPUT125), .A3(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n330_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT126), .B(G197gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1352gat));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n643_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n569_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT63), .B(G211gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n885_), .B2(new_n888_), .ZN(G1354gat));
  INV_X1    g688(.A(G218gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n879_), .B2(new_n609_), .ZN(new_n891_));
  AOI211_X1 g690(.A(G218gat), .B(new_n552_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT127), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n879_), .A2(new_n890_), .A3(new_n577_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n554_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n894_), .B(new_n895_), .C1(new_n890_), .C2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n897_), .ZN(G1355gat));
endmodule


