//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(G50gat), .ZN(new_n205_));
  INV_X1    g004(.A(G29gat), .ZN(new_n206_));
  INV_X1    g005(.A(G36gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT74), .ZN(new_n211_));
  INV_X1    g010(.A(G43gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n213_), .A3(new_n209_), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n212_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n205_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n211_), .A2(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G43gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(G50gat), .A3(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n217_), .A2(new_n221_), .A3(KEYINPUT15), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT15), .B1(new_n217_), .B2(new_n221_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT9), .A3(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT10), .B(G99gat), .Z(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT64), .A3(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n229_), .A2(KEYINPUT9), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT10), .B(G99gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n237_), .B2(G106gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n231_), .A2(new_n234_), .A3(new_n235_), .A4(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT8), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n225_), .B2(new_n226_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G99gat), .A2(G106gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT6), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  NAND3_X1  g044(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n233_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT7), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n248_), .A2(new_n252_), .A3(new_n249_), .A4(new_n233_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n241_), .A2(new_n247_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n228_), .A2(new_n229_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n240_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n240_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n251_), .A2(new_n253_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n227_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n239_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT70), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n239_), .B(new_n262_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n224_), .A2(new_n264_), .A3(KEYINPUT75), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n241_), .A2(new_n247_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n253_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n255_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT8), .ZN(new_n269_));
  INV_X1    g068(.A(new_n227_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n240_), .B(new_n255_), .C1(new_n267_), .C2(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n231_), .A2(new_n238_), .A3(new_n234_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n269_), .A2(new_n271_), .B1(new_n272_), .B2(new_n235_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n217_), .A2(new_n221_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n265_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT75), .B1(new_n224_), .B2(new_n264_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n204_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G190gat), .B(G218gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G134gat), .ZN(new_n280_));
  INV_X1    g079(.A(G162gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT36), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n224_), .A2(new_n264_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n204_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n275_), .A3(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n278_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n282_), .B(KEYINPUT36), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT76), .Z(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n278_), .B2(new_n288_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT37), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n289_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n288_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n285_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n265_), .A3(new_n275_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n298_), .B2(new_n204_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n290_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT77), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n284_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n278_), .A2(new_n288_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n290_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n294_), .B1(new_n306_), .B2(new_n293_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G155gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G183gat), .B(G211gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT17), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT11), .ZN(new_n315_));
  INV_X1    g114(.A(G71gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT67), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G71gat), .ZN(new_n319_));
  INV_X1    g118(.A(G78gat), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n315_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G78gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT11), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G57gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT68), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G57gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G64gat), .ZN(new_n333_));
  INV_X1    g132(.A(G64gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n323_), .A2(new_n327_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n321_), .A2(new_n322_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n338_), .A2(KEYINPUT11), .A3(new_n333_), .A4(new_n335_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(KEYINPUT69), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT69), .B1(new_n337_), .B2(new_n339_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G15gat), .B(G22gat), .ZN(new_n344_));
  INV_X1    g143(.A(G1gat), .ZN(new_n345_));
  INV_X1    g144(.A(G8gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT14), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G1gat), .B(G8gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(G231gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT78), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n350_), .B(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n314_), .B1(new_n343_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n343_), .B2(new_n353_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n313_), .B2(new_n312_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT80), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n337_), .A2(new_n339_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n353_), .B(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n359_), .A2(new_n314_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G120gat), .B(G148gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT5), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G176gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n364_), .B(G204gat), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n337_), .A2(new_n339_), .A3(KEYINPUT12), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n264_), .B2(new_n369_), .ZN(new_n370_));
  AOI211_X1 g169(.A(KEYINPUT71), .B(new_n368_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n341_), .A2(new_n342_), .A3(new_n260_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G230gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n373_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n358_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n273_), .A2(new_n379_), .A3(new_n340_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(KEYINPUT72), .A3(new_n375_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT12), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n343_), .B2(new_n273_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n372_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n343_), .A2(new_n273_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n376_), .B1(new_n386_), .B2(new_n374_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n366_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n366_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n390_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n388_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT13), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n307_), .A2(new_n361_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT81), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n274_), .A2(new_n350_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n350_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n224_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G229gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT84), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n274_), .A2(new_n350_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT83), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n411_), .A2(new_n403_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n412_), .B2(new_n406_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G113gat), .B(G141gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT86), .ZN(new_n415_));
  INV_X1    g214(.A(G169gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G197gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT85), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n413_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT102), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G197gat), .B(G204gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT21), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G211gat), .B(G218gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT21), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT97), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n426_), .A2(new_n432_), .A3(new_n427_), .A4(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n427_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT23), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT89), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT23), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(G183gat), .A3(G190gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(KEYINPUT89), .A3(KEYINPUT23), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT100), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G169gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G176gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G169gat), .A2(G176gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT100), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n445_), .A2(new_n456_), .A3(new_n447_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n449_), .A2(new_n454_), .A3(new_n455_), .A4(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G183gat), .ZN(new_n460_));
  INV_X1    g259(.A(G183gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT25), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT26), .B(G190gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(new_n464_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G169gat), .A2(G176gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT24), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n455_), .A2(KEYINPUT24), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT98), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n465_), .B(new_n468_), .C1(new_n470_), .C2(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n458_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n437_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n435_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT90), .B(G169gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n446_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n469_), .A2(new_n466_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n445_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n459_), .A2(KEYINPUT87), .A3(G183gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n460_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G190gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT26), .ZN(new_n487_));
  AND4_X1   g286(.A1(new_n482_), .A2(new_n484_), .A3(new_n487_), .A4(new_n462_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n486_), .A2(KEYINPUT26), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n488_), .A2(new_n489_), .B1(new_n467_), .B2(new_n466_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n479_), .B1(new_n481_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n474_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n473_), .A2(KEYINPUT20), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G226gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT19), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT20), .B(new_n496_), .C1(new_n474_), .C2(new_n491_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n474_), .A2(new_n458_), .A3(new_n471_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n493_), .A2(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G64gat), .B(G92gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  OAI21_X1  g304(.A(new_n422_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n505_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n437_), .B2(new_n472_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n496_), .B1(new_n510_), .B2(new_n492_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n499_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(new_n497_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT102), .B(new_n508_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n506_), .A2(new_n507_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G225gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G141gat), .ZN(new_n518_));
  INV_X1    g317(.A(G148gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G141gat), .A2(G148gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G155gat), .A2(G162gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G155gat), .A2(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT1), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n520_), .B(new_n521_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n527_));
  OR3_X1    g326(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT2), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n521_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n522_), .B(KEYINPUT93), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(G127gat), .A2(G134gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G127gat), .A2(G134gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(G113gat), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT92), .ZN(new_n545_));
  INV_X1    g344(.A(G113gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n540_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(G120gat), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(G120gat), .B1(new_n543_), .B2(new_n547_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n536_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n536_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n543_), .A2(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(G120gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n555_), .A3(new_n548_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT103), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n549_), .A2(new_n550_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(KEYINPUT103), .A3(new_n552_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n517_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(KEYINPUT4), .A3(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT4), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n551_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n516_), .B(KEYINPUT104), .Z(new_n566_));
  AOI21_X1  g365(.A(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G1gat), .B(G29gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(G85gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT0), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n328_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n517_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n558_), .A2(new_n560_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n574_), .A2(new_n566_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n573_), .A2(new_n575_), .A3(new_n571_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n567_), .A2(KEYINPUT33), .A3(new_n571_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n515_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT105), .ZN(new_n581_));
  INV_X1    g380(.A(new_n571_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n565_), .A2(new_n566_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT107), .B(new_n582_), .C1(new_n583_), .C2(new_n561_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT107), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n572_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(KEYINPUT106), .A2(KEYINPUT20), .ZN(new_n588_));
  OR2_X1    g387(.A1(KEYINPUT106), .A2(KEYINPUT20), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n588_), .B(new_n589_), .C1(new_n474_), .C2(new_n491_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n495_), .B1(new_n512_), .B2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n495_), .B2(new_n493_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n505_), .A2(KEYINPUT32), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n511_), .A2(new_n513_), .A3(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT105), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n515_), .A2(new_n578_), .A3(new_n597_), .A4(new_n579_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n581_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n559_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n600_), .A2(new_n602_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G71gat), .B(G99gat), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n491_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G15gat), .B(G43gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT31), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G227gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n609_), .B(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n606_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n608_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n608_), .B2(new_n615_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n474_), .B1(KEYINPUT29), .B2(new_n536_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT28), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G22gat), .B(G50gat), .Z(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT94), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n622_), .B(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n536_), .A2(KEYINPUT29), .ZN(new_n626_));
  INV_X1    g425(.A(G233gat), .ZN(new_n627_));
  OR2_X1    g426(.A1(KEYINPUT95), .A2(G228gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(KEYINPUT95), .A2(G228gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n626_), .B(new_n630_), .Z(new_n631_));
  XOR2_X1   g430(.A(G78gat), .B(G106gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n625_), .A2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n622_), .A2(new_n624_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n622_), .A2(new_n624_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n633_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n599_), .A2(new_n619_), .A3(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n515_), .A2(KEYINPUT27), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n592_), .A2(new_n508_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n643_), .A2(KEYINPUT108), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(KEYINPUT108), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n644_), .A2(KEYINPUT27), .A3(new_n507_), .A4(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n587_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n619_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n618_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n649_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n421_), .B1(new_n641_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n400_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT109), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT109), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n400_), .A2(new_n657_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G1gat), .A3(new_n649_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT38), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n654_), .A2(new_n398_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n361_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n306_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G1gat), .B1(new_n666_), .B2(new_n649_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(KEYINPUT38), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n667_), .A3(new_n668_), .ZN(G1324gat));
  NAND4_X1  g468(.A1(new_n656_), .A2(new_n346_), .A3(new_n647_), .A4(new_n658_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(new_n665_), .A3(new_n647_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(G8gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(G8gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT110), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n670_), .B(new_n677_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n676_), .A2(KEYINPUT40), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT40), .B1(new_n676_), .B2(new_n678_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1325gat));
  OAI21_X1  g480(.A(G15gat), .B1(new_n666_), .B2(new_n619_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT41), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n659_), .A2(G15gat), .A3(new_n619_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1326gat));
  OAI21_X1  g484(.A(G22gat), .B1(new_n666_), .B2(new_n640_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT42), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT42), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n640_), .A2(G22gat), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n687_), .A2(new_n688_), .B1(new_n659_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT111), .ZN(G1327gat));
  NOR2_X1   g490(.A1(new_n361_), .A2(new_n306_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n662_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n206_), .A3(new_n587_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n641_), .A2(new_n653_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n307_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(KEYINPUT43), .A3(new_n696_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(new_n663_), .A3(new_n398_), .A4(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n421_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT44), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(KEYINPUT44), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n703_), .B(KEYINPUT44), .C1(new_n701_), .C2(new_n421_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n649_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n694_), .B1(new_n708_), .B2(new_n206_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n707_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n207_), .B1(new_n711_), .B2(new_n647_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n693_), .A2(new_n207_), .A3(new_n647_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n714_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n710_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n715_), .A2(new_n716_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n648_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n719_), .B(KEYINPUT46), .C1(new_n207_), .C2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n693_), .A2(new_n212_), .A3(new_n618_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n619_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n212_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT47), .B(new_n723_), .C1(new_n724_), .C2(new_n212_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1330gat));
  NAND3_X1  g528(.A1(new_n693_), .A2(new_n205_), .A3(new_n639_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n640_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n205_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n398_), .A2(new_n420_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n695_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n665_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n328_), .A3(new_n649_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n307_), .A2(new_n361_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n587_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n328_), .B2(new_n740_), .ZN(G1332gat));
  OAI21_X1  g540(.A(G64gat), .B1(new_n735_), .B2(new_n648_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n334_), .A3(new_n647_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n735_), .B2(new_n619_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT49), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n739_), .A2(new_n316_), .A3(new_n618_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n735_), .B2(new_n640_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n739_), .A2(new_n320_), .A3(new_n639_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1335gat));
  NAND2_X1  g553(.A1(new_n734_), .A2(new_n692_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n587_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n699_), .A2(new_n663_), .A3(new_n700_), .A4(new_n733_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n587_), .A2(G85gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1336gat));
  AOI21_X1  g560(.A(G92gat), .B1(new_n756_), .B2(new_n647_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n647_), .A2(G92gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n759_), .B2(new_n763_), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n758_), .B2(new_n619_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n756_), .A2(new_n232_), .A3(new_n618_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT114), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n767_), .B(new_n769_), .ZN(G1338gat));
  OAI21_X1  g569(.A(G106gat), .B1(new_n758_), .B2(new_n640_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT115), .B(G106gat), .C1(new_n758_), .C2(new_n640_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(KEYINPUT52), .A3(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n756_), .A2(new_n233_), .A3(new_n639_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(new_n772_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n775_), .A2(new_n780_), .A3(new_n776_), .A4(new_n778_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1339gat));
  NAND4_X1  g583(.A1(new_n737_), .A2(KEYINPUT117), .A3(new_n421_), .A4(new_n398_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n399_), .B2(new_n420_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(KEYINPUT54), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n786_), .B(new_n789_), .C1(new_n399_), .C2(new_n420_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n269_), .A2(new_n271_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n262_), .B1(new_n794_), .B2(new_n239_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n263_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n369_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT71), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n264_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n384_), .A3(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n380_), .A2(KEYINPUT72), .A3(new_n375_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT72), .B1(new_n380_), .B2(new_n375_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n793_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n798_), .A2(new_n380_), .A3(new_n384_), .A4(new_n799_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n376_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n372_), .A2(new_n382_), .A3(KEYINPUT55), .A4(new_n384_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n365_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n408_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n412_), .B2(new_n408_), .ZN(new_n812_));
  MUX2_X1   g611(.A(new_n812_), .B(new_n413_), .S(new_n418_), .Z(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n808_), .A2(new_n814_), .A3(new_n365_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n810_), .A2(new_n813_), .A3(new_n390_), .A4(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n792_), .B1(new_n816_), .B2(KEYINPUT118), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n696_), .A3(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n810_), .A2(new_n420_), .A3(new_n390_), .A4(new_n815_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n813_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n306_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n664_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n826_), .A2(KEYINPUT57), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n828_), .A3(KEYINPUT57), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n820_), .A2(new_n825_), .A3(new_n827_), .A4(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n791_), .B1(new_n663_), .B2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n647_), .A2(new_n649_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n831_), .A2(new_n651_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834_), .B2(new_n420_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n834_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n838_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n421_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n835_), .B1(new_n841_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g641(.A(new_n554_), .B1(new_n398_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n834_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n554_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n398_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n554_), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n834_), .B2(new_n361_), .ZN(new_n847_));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n361_), .B2(KEYINPUT121), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(KEYINPUT121), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n850_), .B2(new_n851_), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n834_), .B2(new_n664_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n839_), .A2(new_n840_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n696_), .A2(G134gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT122), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n854_), .B2(new_n856_), .ZN(G1343gat));
  INV_X1    g656(.A(new_n650_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n826_), .A2(KEYINPUT57), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n816_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n817_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n861_), .B2(new_n696_), .ZN(new_n862_));
  AND4_X1   g661(.A1(new_n828_), .A2(new_n823_), .A3(KEYINPUT57), .A4(new_n306_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n828_), .B1(new_n826_), .B2(KEYINPUT57), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n361_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n858_), .B(new_n832_), .C1(new_n866_), .C2(new_n791_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT124), .B1(new_n867_), .B2(new_n421_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n830_), .A2(new_n663_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n791_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n650_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n420_), .A4(new_n832_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(new_n869_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n869_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n518_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n868_), .A2(new_n874_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT123), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(G141gat), .A3(new_n875_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n867_), .A2(new_n398_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n519_), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n867_), .A2(new_n663_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT61), .B(G155gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  NOR3_X1   g686(.A1(new_n867_), .A2(new_n281_), .A3(new_n307_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n872_), .A2(new_n664_), .A3(new_n832_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n281_), .B2(new_n889_), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n831_), .A2(new_n651_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n648_), .A2(new_n587_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n891_), .A2(new_n420_), .A3(new_n452_), .A4(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n892_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n421_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n895_), .B2(new_n416_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT62), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n895_), .B2(new_n416_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1348gat));
  NOR2_X1   g699(.A1(new_n894_), .A2(new_n398_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n453_), .ZN(G1349gat));
  INV_X1    g701(.A(new_n463_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n891_), .A2(new_n361_), .A3(new_n903_), .A4(new_n892_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n461_), .B1(new_n894_), .B2(new_n663_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n905_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n894_), .B2(new_n307_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n664_), .A2(new_n464_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n894_), .B2(new_n911_), .ZN(G1351gat));
  OAI211_X1 g711(.A(new_n858_), .B(new_n892_), .C1(new_n866_), .C2(new_n791_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n870_), .A2(new_n871_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n916_), .A2(KEYINPUT126), .A3(new_n858_), .A4(new_n892_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n420_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g719(.A(new_n398_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n918_), .B2(new_n361_), .ZN(new_n924_));
  XOR2_X1   g723(.A(KEYINPUT63), .B(G211gat), .Z(new_n925_));
  AOI211_X1 g724(.A(new_n663_), .B(new_n925_), .C1(new_n915_), .C2(new_n917_), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT127), .B1(new_n924_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n925_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n918_), .A2(new_n361_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n663_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n929_), .B(new_n930_), .C1(new_n931_), .C2(new_n923_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n927_), .A2(new_n932_), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n918_), .B2(new_n664_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n307_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(G218gat), .B2(new_n935_), .ZN(G1355gat));
endmodule


