//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT70), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT64), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n207_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(KEYINPUT9), .A2(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n214_), .B(new_n218_), .C1(KEYINPUT9), .C2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n222_), .B(new_n217_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n224_), .B(new_n225_), .C1(G99gat), .C2(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n221_), .B(new_n227_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n215_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n228_), .B2(new_n215_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(G29gat), .A2(G36gat), .ZN(new_n233_));
  INV_X1    g032(.A(G43gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G29gat), .A2(G36gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G50gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n234_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G43gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(G50gat), .B1(new_n242_), .B2(new_n236_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n238_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(G50gat), .A3(new_n236_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n244_), .A2(KEYINPUT15), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT15), .B1(new_n244_), .B2(new_n248_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n205_), .B(new_n232_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n227_), .A2(new_n221_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n215_), .B1(new_n213_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT8), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n228_), .A2(new_n229_), .A3(new_n215_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n240_), .A2(new_n243_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n220_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT15), .ZN(new_n260_));
  INV_X1    g059(.A(new_n248_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n246_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n244_), .A2(KEYINPUT15), .A3(new_n248_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n205_), .B1(new_n265_), .B2(new_n232_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n204_), .B1(new_n259_), .B2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n232_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n204_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n258_), .A3(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G190gat), .B(G218gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G134gat), .ZN(new_n274_));
  INV_X1    g073(.A(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n267_), .A2(new_n268_), .A3(new_n272_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(new_n272_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n276_), .B(KEYINPUT36), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT72), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n282_));
  AOI211_X1 g081(.A(new_n282_), .B(new_n279_), .C1(new_n267_), .C2(new_n272_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n277_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT104), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT104), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n286_), .B(new_n277_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n291_));
  OAI21_X1  g090(.A(G169gat), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT22), .ZN(new_n297_));
  OAI211_X1 g096(.A(KEYINPUT78), .B(G169gat), .C1(new_n290_), .C2(new_n291_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT76), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT23), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(KEYINPUT23), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G183gat), .ZN(new_n314_));
  INV_X1    g113(.A(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n299_), .A2(KEYINPUT79), .A3(new_n300_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n303_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n296_), .A2(new_n295_), .A3(KEYINPUT75), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(G169gat), .B2(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n310_), .A2(new_n304_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT25), .B(G183gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT24), .B1(new_n320_), .B2(new_n322_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n325_), .A2(new_n327_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334_));
  INV_X1    g133(.A(G204gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT21), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT86), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n338_), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n339_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n334_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n335_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G197gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(G204gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT87), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT21), .ZN(new_n351_));
  OAI21_X1  g150(.A(G204gat), .B1(new_n336_), .B2(new_n337_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n334_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n344_), .A2(new_n355_), .B1(new_n357_), .B2(KEYINPUT21), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n319_), .A2(new_n333_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n300_), .A2(new_n361_), .A3(KEYINPUT24), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n300_), .B2(KEYINPUT24), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n323_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n330_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT94), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n313_), .A2(new_n332_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n312_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT94), .B1(new_n370_), .B2(new_n331_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n363_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n300_), .A2(new_n361_), .A3(KEYINPUT24), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT93), .B(new_n330_), .C1(new_n374_), .C2(new_n323_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n366_), .A2(new_n368_), .A3(new_n371_), .A4(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n300_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G169gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n295_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n327_), .A2(new_n316_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n380_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n342_), .A2(new_n343_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n357_), .A2(KEYINPUT21), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n359_), .A2(new_n390_), .A3(KEYINPUT20), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT19), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT91), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n376_), .A2(new_n387_), .A3(new_n388_), .A4(new_n384_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n393_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n397_), .A2(KEYINPUT20), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n319_), .A2(new_n333_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n389_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT18), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G64gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(G92gat), .Z(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n407_));
  AND4_X1   g206(.A1(KEYINPUT20), .A2(new_n359_), .A3(new_n394_), .A4(new_n390_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n397_), .A2(KEYINPUT20), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT100), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n397_), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n401_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n413_), .B2(new_n393_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT27), .B(new_n407_), .C1(new_n414_), .C2(new_n406_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT27), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n395_), .A2(new_n391_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n406_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n396_), .A2(new_n402_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n406_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT96), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n423_), .A3(new_n407_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n416_), .B1(new_n417_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT1), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(G155gat), .B2(G162gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(G155gat), .A3(G162gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT1), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n434_), .A3(KEYINPUT83), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n437_), .B(KEYINPUT3), .Z(new_n441_));
  XOR2_X1   g240(.A(new_n439_), .B(KEYINPUT2), .Z(new_n442_));
  OAI211_X1 g241(.A(new_n433_), .B(new_n432_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G127gat), .B(G134gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G113gat), .B(G120gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n447_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT82), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n445_), .A2(new_n447_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT97), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n444_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n445_), .A2(new_n447_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n458_), .B2(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n449_), .A2(KEYINPUT82), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n449_), .A2(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n440_), .A2(new_n443_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n457_), .B(KEYINPUT4), .C1(new_n462_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n444_), .A2(new_n455_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n456_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT98), .B(G85gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT0), .B(G57gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n468_), .A2(new_n464_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(new_n472_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n471_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n478_), .B1(new_n484_), .B2(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT29), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n440_), .A2(new_n443_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT28), .ZN(new_n490_));
  INV_X1    g289(.A(G22gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n440_), .A2(new_n443_), .A3(new_n492_), .A4(new_n488_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n238_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G22gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(G50gat), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n444_), .A2(KEYINPUT29), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n389_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n389_), .A2(KEYINPUT84), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G228gat), .A2(G233gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n505_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n389_), .B(new_n502_), .C1(KEYINPUT84), .C2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G78gat), .B(G106gat), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n501_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n501_), .B(KEYINPUT88), .C1(new_n511_), .C2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n451_), .A2(new_n454_), .A3(KEYINPUT31), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n400_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n400_), .A2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n523_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n522_), .B(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n400_), .A2(new_n525_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n526_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G15gat), .B(G43gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G71gat), .B(G99gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n529_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n387_), .A2(new_n388_), .B1(new_n444_), .B2(KEYINPUT29), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n540_), .A2(new_n542_), .A3(new_n507_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n508_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n509_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n512_), .A2(KEYINPUT90), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n501_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n506_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n517_), .A2(new_n539_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n539_), .B1(new_n517_), .B2(new_n553_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n425_), .B(new_n487_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n479_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n471_), .B2(new_n480_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n420_), .A2(new_n423_), .A3(new_n407_), .A4(new_n558_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n484_), .A2(new_n478_), .A3(new_n481_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT33), .B1(new_n560_), .B2(KEYINPUT99), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT33), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n483_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n486_), .B1(new_n414_), .B2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n419_), .A2(new_n566_), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n559_), .A2(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n539_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n515_), .A2(new_n516_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n289_), .B1(new_n556_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G230gat), .ZN(new_n574_));
  INV_X1    g373(.A(G233gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G71gat), .B(G78gat), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT11), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(KEYINPUT11), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(KEYINPUT11), .A3(new_n580_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n220_), .B(new_n586_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT12), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n256_), .B2(new_n220_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n232_), .A2(new_n591_), .A3(new_n585_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n577_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n589_), .A2(KEYINPUT66), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT66), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n587_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n595_), .B(new_n576_), .C1(new_n589_), .C2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n594_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT68), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n594_), .A2(new_n598_), .A3(KEYINPUT68), .A4(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n598_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n232_), .A2(new_n585_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT12), .A3(new_n587_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n576_), .B1(new_n612_), .B2(new_n592_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n603_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT13), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G15gat), .B(G22gat), .ZN(new_n618_));
  INV_X1    g417(.A(G1gat), .ZN(new_n619_));
  INV_X1    g418(.A(G8gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT14), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G1gat), .B(G8gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n265_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n257_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n257_), .B(new_n624_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(new_n296_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(G197gat), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT74), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n637_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n617_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G231gat), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n575_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT16), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(G183gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G211gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n647_), .B(new_n314_), .ZN(new_n650_));
  INV_X1    g449(.A(G211gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n645_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(KEYINPUT73), .A3(new_n627_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n627_), .B1(new_n653_), .B2(KEYINPUT73), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n644_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n644_), .A3(new_n656_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n586_), .A3(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n655_), .A2(new_n644_), .A3(new_n656_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n585_), .B1(new_n661_), .B2(new_n657_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n649_), .A2(new_n652_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(KEYINPUT17), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n662_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n573_), .A2(new_n642_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n667_), .B2(new_n487_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n424_), .A2(new_n417_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n487_), .A3(new_n415_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n517_), .A2(new_n553_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n570_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n571_), .A2(new_n539_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n640_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT101), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n556_), .A2(new_n572_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n640_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n278_), .A2(new_n280_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(KEYINPUT37), .A3(new_n277_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT37), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n284_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n666_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n677_), .A2(new_n680_), .A3(new_n616_), .A4(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(G1gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n486_), .B(KEYINPUT102), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n689_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n690_), .B1(new_n689_), .B2(new_n692_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n668_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT105), .ZN(G1324gat));
  INV_X1    g495(.A(new_n688_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n425_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n620_), .A3(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G8gat), .B1(new_n667_), .B2(new_n425_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT39), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT39), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g503(.A(G15gat), .B1(new_n667_), .B2(new_n570_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT41), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n688_), .A2(G15gat), .A3(new_n570_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1326gat));
  OAI21_X1  g507(.A(G22gat), .B1(new_n667_), .B2(new_n571_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n491_), .A3(new_n671_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1327gat));
  NAND2_X1  g512(.A1(new_n284_), .A2(new_n684_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n682_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT43), .B1(new_n678_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n717_), .B(new_n685_), .C1(new_n556_), .C2(new_n572_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n666_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n721_));
  NAND4_X1  g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n642_), .A4(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n715_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n717_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT43), .B(new_n715_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n720_), .A3(new_n642_), .A4(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(KEYINPUT107), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n692_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G29gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n288_), .A2(new_n666_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n677_), .A2(new_n680_), .A3(new_n616_), .A4(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n487_), .A2(G29gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n734_), .A2(G36gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT45), .B1(new_n739_), .B2(new_n698_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741_));
  NOR4_X1   g540(.A1(new_n734_), .A2(new_n741_), .A3(G36gat), .A4(new_n425_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n722_), .A2(new_n698_), .A3(new_n730_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G36gat), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n737_), .B(new_n738_), .C1(new_n743_), .C2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n739_), .A2(new_n698_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n741_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n742_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT46), .B1(new_n750_), .B2(KEYINPUT108), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n746_), .A2(new_n751_), .ZN(G1329gat));
  NAND4_X1  g551(.A1(new_n722_), .A2(new_n730_), .A3(G43gat), .A4(new_n539_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n234_), .B1(new_n734_), .B2(new_n570_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g555(.A1(new_n722_), .A2(new_n671_), .A3(new_n730_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n671_), .A2(new_n238_), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n757_), .A2(new_n238_), .B1(new_n734_), .B2(new_n758_), .ZN(G1331gat));
  NOR2_X1   g558(.A1(new_n616_), .A2(new_n640_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n678_), .A2(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(new_n687_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n692_), .ZN(new_n763_));
  AND4_X1   g562(.A1(new_n666_), .A2(new_n573_), .A3(new_n641_), .A4(new_n617_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n486_), .A2(G57gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n764_), .B2(new_n698_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT48), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n762_), .A2(new_n767_), .A3(new_n698_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n764_), .B2(new_n539_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT49), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n772_), .A3(new_n539_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  INV_X1    g575(.A(G78gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n764_), .B2(new_n671_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT50), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n762_), .A2(new_n777_), .A3(new_n671_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1335gat));
  NAND2_X1  g580(.A1(new_n761_), .A2(new_n733_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT109), .ZN(new_n783_));
  AOI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n692_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n719_), .A2(new_n720_), .A3(new_n760_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n786_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n487_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n784_), .B1(new_n789_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g589(.A(G92gat), .B1(new_n783_), .B2(new_n698_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n425_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g592(.A1(new_n783_), .A2(new_n216_), .A3(new_n539_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G99gat), .B1(new_n785_), .B2(new_n570_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n783_), .A2(new_n217_), .A3(new_n671_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n719_), .A2(new_n720_), .A3(new_n671_), .A4(new_n760_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(G106gat), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n799_), .B2(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n798_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n698_), .A2(new_n691_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n612_), .B2(new_n592_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n576_), .A2(KEYINPUT112), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n612_), .A2(new_n592_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n577_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n603_), .B(new_n810_), .C1(new_n813_), .C2(new_n808_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n625_), .A2(new_n628_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(G229gat), .A3(G233gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n630_), .A2(new_n626_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n635_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n629_), .A2(new_n635_), .A3(new_n631_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n812_), .A2(KEYINPUT55), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n613_), .B2(new_n811_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n603_), .A4(new_n810_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n815_), .A2(new_n609_), .A3(new_n821_), .A4(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n715_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT115), .B(new_n715_), .C1(new_n828_), .C2(new_n830_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n826_), .A2(new_n829_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT116), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n615_), .A2(new_n821_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n815_), .A2(new_n609_), .A3(new_n640_), .A4(new_n825_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n288_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n838_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT113), .B(KEYINPUT57), .C1(new_n288_), .C2(new_n841_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n666_), .B1(new_n837_), .B2(new_n846_), .ZN(new_n847_));
  AND4_X1   g646(.A1(KEYINPUT111), .A2(new_n666_), .A3(new_n639_), .A4(new_n638_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT111), .B1(new_n666_), .B2(new_n641_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n616_), .B(new_n685_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n554_), .B(new_n806_), .C1(new_n847_), .C2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n640_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n837_), .A2(new_n846_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n720_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n852_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(KEYINPUT117), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n859_), .A2(new_n554_), .A3(new_n806_), .A4(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n853_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n640_), .A2(G113gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT118), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n855_), .B1(new_n865_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n616_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n854_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n616_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n854_), .B2(new_n666_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n720_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G127gat), .ZN(G1342gat));
  NAND2_X1  g675(.A1(new_n715_), .A2(G134gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT119), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n853_), .A2(new_n863_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n861_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n853_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n853_), .B2(new_n288_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(KEYINPUT120), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886_));
  INV_X1    g685(.A(new_n878_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n884_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n886_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n890_), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n806_), .A2(new_n555_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT121), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n640_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n617_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n666_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n894_), .B2(new_n289_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n685_), .A2(new_n275_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n894_), .B2(new_n903_), .ZN(G1347gat));
  AOI21_X1  g703(.A(new_n673_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n425_), .A2(new_n692_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n640_), .A4(new_n907_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n554_), .B(new_n907_), .C1(new_n847_), .C2(new_n852_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT122), .B1(new_n909_), .B2(new_n641_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(G169gat), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n905_), .A2(new_n378_), .A3(new_n640_), .A4(new_n907_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n908_), .A2(new_n910_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  OAI22_X1  g715(.A1(new_n909_), .A2(new_n616_), .B1(KEYINPUT123), .B2(new_n295_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n295_), .A2(KEYINPUT123), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT124), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n917_), .B(new_n919_), .ZN(G1349gat));
  NOR2_X1   g719(.A1(new_n909_), .A2(new_n720_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n328_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n314_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n909_), .B2(new_n685_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n289_), .A2(new_n329_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT125), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n909_), .B2(new_n926_), .ZN(G1351gat));
  AOI21_X1  g726(.A(new_n672_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n425_), .A2(new_n486_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n641_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n348_), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n335_), .A2(KEYINPUT126), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n335_), .A2(KEYINPUT126), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n930_), .A2(new_n616_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n930_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n617_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n937_), .B2(new_n933_), .ZN(G1353gat));
  XOR2_X1   g737(.A(KEYINPUT63), .B(G211gat), .Z(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(new_n666_), .A3(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n930_), .B2(new_n720_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n936_), .B2(new_n289_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n715_), .A2(G218gat), .ZN(new_n945_));
  XOR2_X1   g744(.A(new_n945_), .B(KEYINPUT127), .Z(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n936_), .B2(new_n946_), .ZN(G1355gat));
endmodule


