//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_;
  INV_X1    g000(.A(G228gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n207_), .A2(KEYINPUT3), .B1(new_n209_), .B2(KEYINPUT2), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n208_), .B(new_n211_), .ZN(new_n212_));
  OAI221_X1 g011(.A(new_n210_), .B1(KEYINPUT3), .B2(new_n207_), .C1(new_n212_), .C2(KEYINPUT2), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT91), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G155gat), .B2(G162gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n212_), .A2(new_n206_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT1), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT92), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n216_), .A2(new_n221_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT92), .B1(new_n225_), .B2(new_n219_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n218_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT21), .ZN(new_n230_));
  INV_X1    g029(.A(G204gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G197gat), .ZN(new_n232_));
  INV_X1    g031(.A(G197gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G204gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT93), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n232_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(KEYINPUT94), .B2(new_n232_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n236_), .B(new_n237_), .C1(KEYINPUT21), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n237_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(KEYINPUT21), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n205_), .B1(new_n229_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n222_), .A2(new_n223_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n225_), .A2(KEYINPUT92), .A3(new_n219_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n247_), .A2(new_n248_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n245_), .B(new_n205_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT96), .B1(new_n246_), .B2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G78gat), .B(G106gat), .Z(new_n254_));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n242_), .A2(new_n244_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n255_), .B(new_n251_), .C1(new_n257_), .C2(new_n205_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n253_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT97), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n254_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n228_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n249_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n204_), .B1(new_n265_), .B2(new_n256_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n255_), .B1(new_n266_), .B2(new_n251_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT97), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n253_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n249_), .A2(new_n250_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT28), .ZN(new_n273_));
  XOR2_X1   g072(.A(G22gat), .B(G50gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n261_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n277_), .B(KEYINPUT97), .C1(new_n259_), .C2(new_n260_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT86), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT81), .B(G183gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(G190gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n280_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT83), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT22), .B(G169gat), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT85), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT85), .B1(new_n294_), .B2(G169gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(G176gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n291_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n281_), .B(KEYINPUT84), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT23), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT81), .B(G183gat), .Z(new_n300_));
  INV_X1    g099(.A(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n299_), .A2(KEYINPUT86), .A3(new_n283_), .A4(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n289_), .A2(new_n297_), .A3(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n300_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT82), .B1(new_n308_), .B2(G190gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(G190gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n307_), .B(new_n309_), .C1(KEYINPUT82), .C2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n281_), .A2(new_n282_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n291_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n304_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT20), .B1(new_n320_), .B2(new_n245_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT100), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n313_), .B1(G183gat), .B2(G190gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n292_), .B(KEYINPUT101), .Z(new_n324_));
  OAI211_X1 g123(.A(new_n323_), .B(new_n315_), .C1(new_n324_), .C2(G176gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n286_), .B1(new_n310_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n314_), .B1(new_n317_), .B2(new_n290_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n245_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT100), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n332_), .B(KEYINPUT20), .C1(new_n320_), .C2(new_n245_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n322_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT99), .Z(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n320_), .A2(new_n245_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(KEYINPUT20), .C1(new_n330_), .C2(new_n245_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(new_n337_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT18), .B(G64gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  AND3_X1   g145(.A1(new_n339_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT102), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G120gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT89), .B(G113gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n227_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n350_), .B1(new_n355_), .B2(KEYINPUT4), .ZN(new_n356_));
  INV_X1    g155(.A(new_n354_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n249_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n358_), .A3(KEYINPUT4), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n227_), .A2(KEYINPUT102), .A3(new_n361_), .A4(new_n354_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n356_), .A2(new_n359_), .A3(new_n360_), .A4(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364_));
  INV_X1    g163(.A(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  AND2_X1   g167(.A1(new_n355_), .A2(new_n358_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n363_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n356_), .A2(new_n359_), .A3(new_n370_), .A4(new_n362_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n360_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n368_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n372_), .B1(new_n378_), .B2(KEYINPUT103), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n376_), .A2(new_n377_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT103), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n381_), .A3(new_n377_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n349_), .A2(new_n379_), .A3(new_n380_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n339_), .A2(KEYINPUT104), .A3(new_n342_), .A4(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n373_), .A2(new_n374_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n368_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n376_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n339_), .A2(new_n342_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n384_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT104), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n341_), .A2(new_n337_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n394_), .B2(new_n390_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n385_), .B(new_n388_), .C1(new_n391_), .C2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n279_), .A2(new_n383_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n346_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(KEYINPUT27), .C1(new_n389_), .C2(new_n400_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n276_), .B(new_n278_), .C1(new_n403_), .C2(new_n388_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G15gat), .B(G43gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G71gat), .B(G99gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n320_), .B(KEYINPUT30), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(KEYINPUT87), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(KEYINPUT87), .B2(new_n410_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n354_), .B(KEYINPUT31), .Z(new_n413_));
  AND2_X1   g212(.A1(new_n413_), .A2(KEYINPUT88), .ZN(new_n414_));
  INV_X1    g213(.A(new_n410_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n409_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n412_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n397_), .A2(new_n404_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT105), .ZN(new_n423_));
  INV_X1    g222(.A(new_n388_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n399_), .A2(new_n402_), .A3(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n423_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n429_));
  NAND2_X1  g228(.A1(G232gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT67), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n435_));
  AND2_X1   g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT7), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT8), .ZN(new_n443_));
  XOR2_X1   g242(.A(G85gat), .B(G92gat), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT68), .B1(new_n437_), .B2(new_n438_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n436_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n432_), .A2(KEYINPUT67), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT68), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n446_), .A2(new_n453_), .A3(new_n441_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n444_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT69), .B1(new_n455_), .B2(KEYINPUT8), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT69), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n457_), .B(new_n443_), .C1(new_n454_), .C2(new_n444_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n445_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G43gat), .B(G50gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(G29gat), .B(G36gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n461_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n465_));
  INV_X1    g264(.A(G92gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n365_), .B2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n467_), .A2(KEYINPUT9), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(KEYINPUT9), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n468_), .B(new_n469_), .C1(G85gat), .C2(G92gat), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n470_), .A2(KEYINPUT66), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT10), .B(G99gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(G106gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT64), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(KEYINPUT66), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n471_), .A2(new_n439_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n459_), .A2(new_n464_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n464_), .B(KEYINPUT15), .Z(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n459_), .B2(new_n476_), .ZN(new_n480_));
  OAI211_X1 g279(.A(KEYINPUT35), .B(new_n431_), .C1(new_n478_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n431_), .A2(KEYINPUT35), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n431_), .A2(KEYINPUT35), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .A4(new_n477_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G190gat), .B(G218gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G134gat), .B(G162gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND4_X1  g289(.A1(new_n481_), .A2(new_n485_), .A3(new_n487_), .A4(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n481_), .A2(new_n485_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n490_), .B(KEYINPUT36), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n492_), .A2(KEYINPUT78), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT78), .B1(new_n492_), .B2(new_n493_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G57gat), .B(G64gat), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G71gat), .B(G78gat), .ZN(new_n503_));
  OR3_X1    g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n503_), .A3(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507_));
  INV_X1    g306(.A(G1gat), .ZN(new_n508_));
  INV_X1    g307(.A(G8gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G8gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n506_), .B(new_n513_), .Z(new_n514_));
  AND2_X1   g313(.A1(G231gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G127gat), .B(G155gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G211gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT16), .B(G183gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(KEYINPUT79), .A3(KEYINPUT17), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n522_), .B1(KEYINPUT17), .B2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n516_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n493_), .B(KEYINPUT77), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n492_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT37), .A3(new_n491_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n498_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n428_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n464_), .B(new_n513_), .Z(new_n532_));
  INV_X1    g331(.A(new_n464_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n513_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n479_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n513_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  MUX2_X1   g336(.A(new_n532_), .B(new_n536_), .S(new_n537_), .Z(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n233_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT80), .B(G169gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n538_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n459_), .A2(new_n476_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n506_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n459_), .A2(new_n476_), .A3(new_n506_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n548_), .A2(KEYINPUT70), .A3(new_n550_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT70), .B1(new_n548_), .B2(new_n550_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n545_), .A2(KEYINPUT12), .A3(new_n546_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n552_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT72), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n552_), .B(new_n566_), .C1(new_n555_), .C2(new_n559_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n560_), .A2(KEYINPUT73), .A3(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n571_), .A2(new_n576_), .A3(new_n577_), .A4(new_n572_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n531_), .A2(new_n544_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n508_), .A3(new_n388_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT38), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n544_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n526_), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n587_), .A2(KEYINPUT106), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n428_), .A2(new_n496_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT106), .B1(new_n587_), .B2(new_n588_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n424_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(G1324gat));
  NAND3_X1  g393(.A1(new_n584_), .A2(new_n509_), .A3(new_n403_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n589_), .A2(new_n591_), .A3(new_n403_), .A4(new_n590_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(G8gat), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n596_), .B2(G8gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g400(.A(G15gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n420_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n584_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n589_), .A2(new_n591_), .A3(new_n603_), .A4(new_n590_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G15gat), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT107), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT41), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(KEYINPUT107), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n604_), .B1(new_n610_), .B2(new_n611_), .ZN(G1326gat));
  INV_X1    g411(.A(G22gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n279_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n584_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n589_), .A2(new_n591_), .A3(new_n614_), .A4(new_n590_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G22gat), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT108), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT42), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(KEYINPUT108), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n615_), .B1(new_n621_), .B2(new_n622_), .ZN(G1327gat));
  NAND3_X1  g422(.A1(new_n583_), .A2(new_n544_), .A3(new_n588_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n496_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n428_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT110), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n624_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n388_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n498_), .A2(new_n529_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT109), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT109), .B1(new_n498_), .B2(new_n529_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n428_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT43), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n428_), .A2(new_n638_), .A3(new_n632_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n624_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT44), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(G29gat), .A3(new_n388_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(KEYINPUT44), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n631_), .B1(new_n642_), .B2(new_n643_), .ZN(G1328gat));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n403_), .A3(new_n643_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n628_), .A2(new_n647_), .A3(new_n403_), .A4(new_n629_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n646_), .A2(KEYINPUT46), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND4_X1  g453(.A1(new_n641_), .A2(G43gat), .A3(new_n603_), .A4(new_n643_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n628_), .A2(new_n603_), .A3(new_n629_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT111), .ZN(new_n657_));
  INV_X1    g456(.A(G43gat), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n630_), .B2(new_n614_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n641_), .A2(G50gat), .A3(new_n643_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n614_), .ZN(G1331gat));
  NOR2_X1   g464(.A1(new_n583_), .A2(new_n544_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n531_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G57gat), .B1(new_n667_), .B2(new_n388_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT112), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n590_), .A2(new_n526_), .A3(new_n666_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(G57gat), .A3(new_n388_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT113), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n670_), .B2(new_n403_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n667_), .A2(new_n675_), .A3(new_n403_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1333gat));
  INV_X1    g478(.A(G71gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n670_), .B2(new_n603_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT49), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n680_), .A3(new_n603_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1334gat));
  INV_X1    g483(.A(G78gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n670_), .B2(new_n614_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT50), .Z(new_n687_));
  NOR2_X1   g486(.A1(new_n279_), .A2(G78gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT114), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n667_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1335gat));
  NAND3_X1  g490(.A1(new_n582_), .A2(new_n543_), .A3(new_n588_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n626_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n388_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n424_), .A2(new_n365_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(G1336gat));
  AOI21_X1  g496(.A(G92gat), .B1(new_n693_), .B2(new_n403_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n403_), .A2(G92gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT115), .Z(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n695_), .B2(new_n700_), .ZN(G1337gat));
  NAND2_X1  g500(.A1(new_n695_), .A2(new_n603_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n420_), .A2(new_n472_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n702_), .A2(G99gat), .B1(new_n693_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT116), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT51), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n704_), .B(new_n706_), .ZN(G1338gat));
  INV_X1    g506(.A(G106gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n695_), .B2(new_n614_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT118), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(KEYINPUT117), .A3(new_n710_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT117), .ZN(new_n713_));
  INV_X1    g512(.A(new_n692_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n632_), .B(new_n633_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n638_), .B1(new_n715_), .B2(new_n428_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n639_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n614_), .B(new_n714_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G106gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n713_), .B1(new_n719_), .B2(KEYINPUT52), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT118), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n721_), .A3(KEYINPUT52), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n711_), .A2(new_n712_), .A3(new_n720_), .A4(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n693_), .A2(new_n708_), .A3(new_n614_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1339gat));
  NOR2_X1   g529(.A1(new_n403_), .A2(new_n424_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n544_), .A2(new_n570_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n548_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n551_), .B1(new_n559_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT12), .B1(new_n545_), .B2(new_n546_), .ZN(new_n738_));
  AOI211_X1 g537(.A(new_n556_), .B(new_n506_), .C1(new_n459_), .C2(new_n476_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(KEYINPUT55), .C1(new_n554_), .C2(new_n553_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n737_), .A3(new_n741_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n742_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT56), .B1(new_n742_), .B2(new_n567_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n733_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n542_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n536_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n537_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n537_), .B2(new_n532_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n538_), .A2(new_n746_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n571_), .A2(new_n572_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n745_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT57), .B1(new_n753_), .B2(new_n496_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n755_), .B(new_n625_), .C1(new_n745_), .C2(new_n752_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n570_), .B(new_n751_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n742_), .A2(new_n567_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n742_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(KEYINPUT58), .A3(new_n570_), .A4(new_n751_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n760_), .A2(new_n766_), .A3(new_n632_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n526_), .B1(new_n757_), .B2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n530_), .A2(new_n581_), .A3(new_n543_), .A4(new_n580_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n422_), .B(new_n731_), .C1(new_n768_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G113gat), .B1(new_n773_), .B2(new_n544_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT59), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n422_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n732_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n752_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n496_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n755_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n753_), .A2(KEYINPUT57), .A3(new_n496_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n767_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n588_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n769_), .A2(KEYINPUT54), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n769_), .A2(KEYINPUT54), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n777_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT59), .A3(new_n731_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n543_), .B1(new_n776_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n774_), .B1(new_n790_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g590(.A(KEYINPUT60), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n583_), .B2(G120gat), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n773_), .B(new_n793_), .C1(new_n792_), .C2(G120gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n583_), .B1(new_n776_), .B2(new_n789_), .ZN(new_n795_));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT120), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n794_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1341gat));
  AOI21_X1  g600(.A(G127gat), .B1(new_n773_), .B2(new_n526_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n776_), .A2(new_n789_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n526_), .A2(G127gat), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT121), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n802_), .B1(new_n803_), .B2(new_n805_), .ZN(G1342gat));
  XOR2_X1   g605(.A(KEYINPUT122), .B(G134gat), .Z(new_n807_));
  AOI22_X1  g606(.A1(new_n783_), .A2(new_n588_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n731_), .ZN(new_n809_));
  NOR4_X1   g608(.A1(new_n808_), .A2(new_n775_), .A3(new_n777_), .A4(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT59), .B1(new_n788_), .B2(new_n731_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n632_), .B(new_n807_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n772_), .B2(new_n496_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n812_), .A2(KEYINPUT123), .A3(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1343gat));
  NOR3_X1   g618(.A1(new_n808_), .A2(new_n279_), .A3(new_n603_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n731_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n544_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n582_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n526_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  AOI21_X1  g627(.A(G162gat), .B1(new_n821_), .B2(new_n625_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n715_), .A2(G162gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n821_), .B2(new_n830_), .ZN(G1347gat));
  NAND2_X1  g630(.A1(new_n403_), .A2(new_n424_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n788_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n544_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(G169gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n836_), .B2(G169gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(KEYINPUT124), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n834_), .A2(KEYINPUT124), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n543_), .A2(new_n324_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n838_), .A2(new_n839_), .B1(new_n843_), .B2(new_n844_), .ZN(G1348gat));
  OAI21_X1  g644(.A(G176gat), .B1(new_n834_), .B2(new_n583_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n583_), .A2(G176gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n843_), .B2(new_n847_), .ZN(G1349gat));
  AOI21_X1  g647(.A(new_n287_), .B1(new_n835_), .B2(new_n526_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n842_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n588_), .B1(new_n850_), .B2(new_n840_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n326_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(G1350gat));
  OAI211_X1 g652(.A(new_n310_), .B(new_n625_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n850_), .A2(new_n840_), .B1(new_n498_), .B2(new_n529_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n301_), .ZN(G1351gat));
  NAND3_X1  g655(.A1(new_n820_), .A2(new_n544_), .A3(new_n833_), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n857_), .A2(KEYINPUT125), .A3(new_n233_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n233_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT125), .B1(new_n857_), .B2(new_n233_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(G1352gat));
  AND2_X1   g660(.A1(new_n820_), .A2(new_n833_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n582_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g663(.A(KEYINPUT63), .B(G211gat), .Z(new_n865_));
  AND3_X1   g664(.A1(new_n862_), .A2(new_n526_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n526_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1354gat));
  AOI21_X1  g668(.A(G218gat), .B1(new_n862_), .B2(new_n625_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n632_), .A2(G218gat), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(KEYINPUT126), .Z(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n862_), .B2(new_n872_), .ZN(G1355gat));
endmodule


