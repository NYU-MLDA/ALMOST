//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT86), .B(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n207_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n215_));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT87), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n219_), .B(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n212_), .B(new_n216_), .C1(new_n225_), .C2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n223_), .A2(KEYINPUT88), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT88), .B1(new_n223_), .B2(new_n228_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n206_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n215_), .A2(KEYINPUT87), .A3(new_n216_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT87), .B1(new_n215_), .B2(new_n216_), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n213_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n222_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n228_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n206_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n231_), .A2(KEYINPUT101), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT101), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n241_), .B(new_n206_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n202_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT103), .B(KEYINPUT4), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n231_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n231_), .A2(KEYINPUT101), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n237_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n247_), .A2(KEYINPUT4), .A3(new_n242_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT102), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n239_), .A2(KEYINPUT102), .A3(KEYINPUT4), .A4(new_n242_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n246_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n244_), .B1(new_n253_), .B2(new_n202_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT0), .B(G57gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G85gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(G1gat), .B(G29gat), .Z(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT106), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n244_), .B(new_n258_), .C1(new_n253_), .C2(new_n202_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n253_), .A2(new_n202_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(KEYINPUT106), .A3(new_n244_), .A4(new_n258_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G36gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT100), .B(G8gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT79), .B(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT80), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G190gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT26), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n274_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(G183gat), .A3(G190gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT82), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n278_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n285_), .A2(KEYINPUT24), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n282_), .A2(new_n287_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n274_), .A2(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G169gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT83), .B1(new_n299_), .B2(KEYINPUT22), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT84), .B(G176gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT22), .B(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n298_), .B(new_n286_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n295_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT92), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT21), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n307_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n311_), .B1(new_n315_), .B2(KEYINPUT21), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n273_), .B1(new_n306_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n278_), .A2(KEYINPUT26), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n280_), .A2(new_n279_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n283_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n297_), .A2(KEYINPUT95), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT95), .B1(new_n297_), .B2(new_n324_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n287_), .B(new_n322_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT96), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n297_), .A2(new_n324_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT95), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n325_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(KEYINPUT96), .A3(new_n287_), .A4(new_n322_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n291_), .A2(new_n278_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n293_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT97), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n302_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n301_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n340_), .A3(new_n286_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n330_), .A2(new_n335_), .A3(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n317_), .B(new_n320_), .C1(new_n316_), .C2(new_n342_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(KEYINPUT98), .A3(new_n316_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT98), .B1(new_n342_), .B2(new_n316_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT20), .B1(new_n306_), .B2(new_n316_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n272_), .B(new_n343_), .C1(new_n347_), .C2(new_n320_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT107), .ZN(new_n349_));
  INV_X1    g148(.A(new_n316_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n341_), .A3(new_n328_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n317_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n319_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n345_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(KEYINPUT98), .A3(new_n316_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n357_), .B2(new_n319_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n272_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n319_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT107), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n272_), .A4(new_n343_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n349_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT27), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n343_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n359_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n348_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n266_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G106gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n373_));
  NAND2_X1  g172(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(G233gat), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n373_), .B1(new_n316_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n236_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n223_), .A2(KEYINPUT88), .A3(new_n228_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n382_), .B2(KEYINPUT29), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n236_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n316_), .B(new_n385_), .C1(new_n387_), .C2(new_n378_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n377_), .ZN(new_n389_));
  AOI221_X4 g188(.A(G78gat), .B1(new_n383_), .B2(KEYINPUT91), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G78gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n383_), .A2(KEYINPUT91), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n372_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n385_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT29), .B1(new_n229_), .B2(new_n230_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n378_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n377_), .B1(new_n399_), .B2(new_n316_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n393_), .ZN(new_n401_));
  OAI21_X1  g200(.A(G78gat), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(G106gat), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n395_), .A2(new_n404_), .A3(KEYINPUT94), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n380_), .A2(new_n386_), .A3(new_n381_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  XNOR2_X1  g207(.A(G22gat), .B(G50gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n395_), .A2(KEYINPUT94), .A3(new_n404_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT94), .B1(new_n395_), .B2(new_n404_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n414_), .B2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n371_), .A2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n272_), .A2(KEYINPUT32), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n358_), .A2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n366_), .A2(new_n417_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n263_), .A2(new_n265_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n239_), .A2(G225gat), .A3(G233gat), .A4(new_n242_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n253_), .A2(KEYINPUT105), .A3(new_n202_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT105), .B1(new_n253_), .B2(new_n202_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n258_), .B(new_n421_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT104), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n260_), .A2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n367_), .A2(new_n348_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n254_), .B(new_n259_), .C1(new_n425_), .C2(KEYINPUT33), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n424_), .A2(new_n427_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT94), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n390_), .A2(new_n394_), .A3(new_n372_), .ZN(new_n432_));
  AOI21_X1  g231(.A(G106gat), .B1(new_n402_), .B2(new_n403_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n410_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n412_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n420_), .A2(new_n430_), .A3(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n306_), .B(KEYINPUT30), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(new_n206_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT85), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n443_), .B(KEYINPUT31), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n441_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n441_), .A2(new_n444_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n441_), .A2(new_n444_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n416_), .A2(new_n439_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT108), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n263_), .A2(new_n265_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n455_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G29gat), .B(G36gat), .ZN(new_n462_));
  INV_X1    g261(.A(G43gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G50gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT77), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n464_), .B(G50gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT77), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G1gat), .B(G8gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(G15gat), .A2(G22gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G15gat), .A2(G22gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G1gat), .A2(G8gat), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n475_), .A2(new_n476_), .B1(KEYINPUT14), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n474_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n471_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n467_), .A2(new_n470_), .A3(new_n479_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n467_), .A2(new_n470_), .A3(KEYINPUT78), .A4(new_n479_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n466_), .B(KEYINPUT15), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n479_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n485_), .A3(new_n481_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(new_n299_), .ZN(new_n494_));
  INV_X1    g293(.A(G197gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n488_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G190gat), .B(G218gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G134gat), .ZN(new_n504_));
  INV_X1    g303(.A(G162gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT36), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT71), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(KEYINPUT71), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  NOR2_X1   g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(KEYINPUT67), .A3(new_n519_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n515_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G85gat), .B(G92gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n512_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(KEYINPUT65), .A3(new_n372_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT65), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT10), .B(G99gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n523_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n525_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT9), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(G85gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(G85gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(KEYINPUT9), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G92gat), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n532_), .A2(new_n533_), .A3(new_n535_), .A4(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(KEYINPUT8), .B(new_n534_), .C1(new_n515_), .C2(new_n520_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n526_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n544_), .A2(KEYINPUT70), .A3(new_n466_), .A4(new_n526_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n543_), .B2(new_n468_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n489_), .A2(new_n543_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT34), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n552_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n554_), .B1(new_n548_), .B2(new_n555_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n510_), .B(new_n511_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n506_), .A4(new_n556_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n502_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n507_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n563_), .B1(new_n502_), .B2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G57gat), .B(G64gat), .Z(new_n568_));
  INV_X1    g367(.A(KEYINPUT11), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(G71gat), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n568_), .A2(new_n569_), .B1(new_n572_), .B2(new_n391_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT68), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n571_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n568_), .A2(new_n569_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n391_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT68), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n570_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n526_), .A3(new_n544_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n543_), .A2(new_n584_), .A3(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT64), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT69), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT69), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n588_), .A2(new_n593_), .A3(new_n590_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n586_), .A2(KEYINPUT12), .A3(new_n587_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n587_), .A2(KEYINPUT12), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n592_), .B(new_n594_), .C1(new_n597_), .C2(new_n590_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G120gat), .B(G148gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G204gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(G176gat), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n598_), .A2(new_n603_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT13), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n598_), .A2(new_n603_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n479_), .B(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(new_n585_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT16), .B(G183gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n585_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n615_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT74), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n614_), .B(new_n585_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n621_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n620_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT75), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(KEYINPUT75), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n624_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n628_), .A2(KEYINPUT75), .ZN(new_n632_));
  INV_X1    g431(.A(new_n624_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(KEYINPUT75), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n631_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n567_), .A2(new_n612_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n501_), .B1(new_n638_), .B2(KEYINPUT76), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n461_), .A2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n638_), .A2(KEYINPUT76), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n642_), .A2(G1gat), .A3(new_n266_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT38), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT109), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT109), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n637_), .A2(new_n566_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n461_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n612_), .A2(new_n501_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n266_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n647_), .B1(new_n653_), .B2(G1gat), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n645_), .B(new_n646_), .C1(new_n654_), .C2(new_n643_), .ZN(G1324gat));
  OR3_X1    g454(.A1(new_n642_), .A2(G8gat), .A3(new_n370_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n370_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n649_), .A2(new_n650_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n658_), .A2(new_n659_), .A3(G8gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n658_), .B2(G8gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n656_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n454_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n651_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT41), .ZN(new_n668_));
  INV_X1    g467(.A(new_n642_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n651_), .A2(new_n415_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G22gat), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(KEYINPUT42), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(KEYINPUT42), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n438_), .A2(G22gat), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT110), .Z(new_n677_));
  OAI22_X1  g476(.A1(new_n674_), .A2(new_n675_), .B1(new_n642_), .B2(new_n677_), .ZN(G1327gat));
  NOR3_X1   g477(.A1(new_n612_), .A2(new_n636_), .A3(new_n501_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n461_), .A2(new_n566_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n652_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n461_), .A2(new_n682_), .A3(new_n567_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n461_), .B2(new_n567_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(G29gat), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n679_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n266_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n681_), .B1(new_n688_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n679_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n460_), .A2(new_n459_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n416_), .A2(new_n439_), .A3(new_n454_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n567_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT43), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n461_), .A2(new_n682_), .A3(new_n567_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n370_), .B1(new_n701_), .B2(KEYINPUT44), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n694_), .B1(new_n702_), .B2(new_n687_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n680_), .A2(new_n694_), .A3(new_n657_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n693_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n701_), .A2(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n689_), .A2(new_n657_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G36gat), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n712_), .ZN(G1329gat));
  NAND3_X1  g512(.A1(new_n461_), .A2(new_n566_), .A3(new_n679_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n463_), .B1(new_n714_), .B2(new_n454_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT111), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n687_), .A2(G43gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n689_), .A2(new_n666_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n721_), .B(new_n716_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n680_), .B2(new_n415_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n708_), .A2(new_n465_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n690_), .A2(new_n438_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n611_), .A2(new_n500_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n649_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(G57gat), .A3(new_n652_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n563_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(KEYINPUT37), .B2(new_n565_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n461_), .A2(new_n636_), .A3(new_n732_), .A4(new_n728_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n266_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(G57gat), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT112), .ZN(G1332gat));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n729_), .A2(new_n657_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n739_), .A3(G64gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n738_), .B2(G64gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n737_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n738_), .A2(G64gat), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT113), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(KEYINPUT48), .A3(new_n740_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n733_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n370_), .A2(G64gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT114), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n743_), .A2(new_n746_), .A3(new_n750_), .ZN(G1333gat));
  NAND2_X1  g550(.A1(new_n649_), .A2(new_n728_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G71gat), .B1(new_n752_), .B2(new_n454_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n572_), .A3(new_n666_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n752_), .B2(new_n438_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n747_), .A2(new_n391_), .A3(new_n415_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n728_), .A2(new_n637_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n461_), .A2(new_n566_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G85gat), .B1(new_n763_), .B2(new_n652_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n266_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n763_), .B2(new_n657_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n657_), .A2(G92gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n765_), .B2(new_n769_), .ZN(G1337gat));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n666_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G99gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n527_), .A3(new_n666_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT51), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n776_), .A3(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n763_), .A2(new_n372_), .A3(new_n415_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n415_), .B(new_n762_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT116), .Z(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n786_), .B(new_n779_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n595_), .A2(new_n590_), .A3(new_n596_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n590_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(KEYINPUT55), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n590_), .B(new_n796_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n603_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(new_n603_), .C1(new_n794_), .C2(new_n797_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n799_), .A2(new_n500_), .A3(new_n608_), .A4(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n490_), .A2(new_n486_), .A3(new_n481_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n496_), .A3(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n499_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n802_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n565_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n799_), .A2(new_n801_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n608_), .A4(new_n806_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n799_), .A2(new_n608_), .A3(new_n806_), .A4(new_n801_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n567_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n811_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n808_), .A2(new_n565_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n812_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n637_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n732_), .A2(new_n611_), .A3(new_n501_), .A4(new_n636_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT54), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n657_), .A2(new_n266_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n457_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n500_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n825_), .A2(new_n826_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(KEYINPUT119), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n457_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(KEYINPUT119), .ZN(new_n834_));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n501_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n829_), .B1(new_n837_), .B2(G113gat), .ZN(G1340gat));
  XOR2_X1   g637(.A(KEYINPUT120), .B(G120gat), .Z(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n611_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n839_), .B2(KEYINPUT60), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n827_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n611_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n839_), .ZN(G1341gat));
  NOR2_X1   g645(.A1(KEYINPUT122), .A2(G127gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(G127gat), .B1(new_n637_), .B2(KEYINPUT122), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI211_X1 g648(.A(new_n847_), .B(new_n849_), .C1(new_n833_), .C2(new_n836_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G127gat), .B1(new_n828_), .B2(new_n636_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT123), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n853_));
  INV_X1    g652(.A(new_n851_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n833_), .A2(new_n836_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n848_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n853_), .B(new_n854_), .C1(new_n856_), .C2(new_n847_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n852_), .A2(new_n857_), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n828_), .B2(new_n566_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n855_), .A2(G134gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n567_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n438_), .A2(new_n666_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n830_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n830_), .A2(KEYINPUT124), .A3(new_n862_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n501_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  AOI21_X1  g668(.A(new_n611_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n870_));
  INV_X1    g669(.A(G148gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n865_), .A2(new_n866_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n873_), .A2(new_n636_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n636_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1346gat));
  AOI21_X1  g676(.A(G162gat), .B1(new_n873_), .B2(new_n566_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n505_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n567_), .B2(new_n879_), .ZN(G1347gat));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n652_), .A2(new_n454_), .A3(new_n370_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n819_), .B1(new_n808_), .B2(new_n565_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n811_), .B(new_n566_), .C1(new_n802_), .C2(new_n807_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n636_), .B1(new_n885_), .B2(new_n818_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n823_), .B(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n438_), .B(new_n882_), .C1(new_n886_), .C2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n881_), .B1(new_n889_), .B2(new_n501_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n415_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n891_), .A2(KEYINPUT125), .A3(new_n500_), .A4(new_n882_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(G169gat), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n889_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n500_), .A3(new_n339_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n890_), .A2(KEYINPUT62), .A3(new_n892_), .A4(G169gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n895_), .A2(KEYINPUT126), .A3(new_n897_), .A4(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1348gat));
  INV_X1    g702(.A(new_n891_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT127), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n905_), .A2(G176gat), .A3(new_n882_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n896_), .A2(new_n612_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n906_), .A2(new_n612_), .B1(new_n301_), .B2(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n889_), .A2(new_n637_), .A3(new_n280_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n636_), .A3(new_n882_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n291_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n889_), .B2(new_n732_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n566_), .A2(new_n279_), .A3(new_n321_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n889_), .B2(new_n913_), .ZN(G1351gat));
  AND2_X1   g713(.A1(new_n825_), .A2(new_n862_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n652_), .A2(new_n370_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n501_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n495_), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n611_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g720(.A1(new_n917_), .A2(new_n637_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT63), .B(G211gat), .Z(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n917_), .A2(new_n926_), .A3(new_n732_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n915_), .A2(new_n566_), .A3(new_n916_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1355gat));
endmodule


