//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT79), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT79), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT24), .B1(new_n202_), .B2(new_n203_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT80), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n207_), .A2(KEYINPUT80), .A3(new_n208_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n211_), .A2(KEYINPUT81), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n207_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n212_), .A2(new_n215_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT81), .B1(new_n223_), .B2(new_n211_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(new_n202_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(new_n219_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(new_n230_), .B2(new_n219_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(KEYINPUT30), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT30), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  INV_X1    g037(.A(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(G15gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n234_), .A2(KEYINPUT82), .A3(new_n237_), .A4(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n234_), .A2(KEYINPUT82), .A3(new_n237_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT82), .B1(new_n234_), .B2(new_n237_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT85), .B(new_n245_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT86), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(new_n245_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT84), .A3(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n260_), .A2(KEYINPUT84), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT31), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n254_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n264_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT90), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(KEYINPUT21), .A3(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n271_), .B(KEYINPUT21), .Z(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT3), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT2), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT87), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n285_), .B1(KEYINPUT1), .B2(new_n283_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(KEYINPUT1), .B2(new_n283_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n277_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n279_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n276_), .B1(new_n292_), .B2(KEYINPUT29), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G228gat), .A2(G233gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n276_), .B2(KEYINPUT89), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n293_), .B(new_n295_), .Z(new_n296_));
  XOR2_X1   g095(.A(G22gat), .B(G50gat), .Z(new_n297_));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n298_), .A3(new_n291_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT88), .ZN(new_n301_));
  INV_X1    g100(.A(new_n291_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n298_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n300_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n297_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G78gat), .B(G106gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT91), .ZN(new_n311_));
  INV_X1    g110(.A(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n304_), .B1(new_n303_), .B2(new_n298_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT88), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n297_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n300_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n308_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n310_), .B1(new_n308_), .B2(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n296_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n306_), .A2(new_n307_), .A3(new_n297_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n315_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n309_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n308_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n296_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT99), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n303_), .B1(new_n262_), .B2(new_n261_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n259_), .A2(new_n260_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n287_), .A2(new_n331_), .A3(new_n291_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT4), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT4), .B1(new_n292_), .B2(new_n263_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT96), .B(G85gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT0), .B(G57gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n292_), .A2(new_n263_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n303_), .A2(new_n331_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n335_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n338_), .A2(new_n344_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n338_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n329_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n338_), .A2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n343_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n338_), .A2(new_n344_), .A3(new_n348_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(KEYINPUT99), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n225_), .A2(new_n276_), .A3(new_n233_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  INV_X1    g157(.A(new_n229_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n227_), .A2(KEYINPUT95), .B1(new_n220_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(KEYINPUT95), .B2(new_n227_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n210_), .A2(new_n220_), .A3(new_n218_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n214_), .B(KEYINPUT94), .ZN(new_n363_));
  INV_X1    g162(.A(new_n213_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n361_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n366_), .B2(new_n275_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n357_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT93), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n366_), .B2(new_n275_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n235_), .B2(new_n275_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n371_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT18), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n368_), .A2(new_n373_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT98), .B1(new_n368_), .B2(new_n373_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT98), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n357_), .A2(new_n391_), .A3(new_n367_), .A4(new_n372_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n376_), .A2(new_n377_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n384_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n389_), .B1(new_n386_), .B2(new_n383_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n388_), .A2(new_n389_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n268_), .A2(new_n328_), .A3(new_n356_), .A4(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n383_), .A2(KEYINPUT32), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n379_), .A2(new_n399_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n400_), .B(new_n401_), .C1(new_n350_), .C2(new_n349_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n345_), .A2(new_n346_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n336_), .B1(new_n403_), .B2(KEYINPUT4), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n347_), .B1(new_n404_), .B2(new_n335_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NOR4_X1   g205(.A1(new_n405_), .A2(KEYINPUT97), .A3(new_n406_), .A4(new_n344_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT97), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n350_), .B2(KEYINPUT33), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n333_), .A2(new_n337_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n334_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n403_), .A2(new_n334_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(new_n343_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n387_), .B(new_n385_), .C1(new_n415_), .C2(new_n350_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n402_), .B1(new_n410_), .B2(new_n416_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n320_), .A2(new_n326_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n417_), .A2(new_n328_), .B1(new_n418_), .B2(new_n397_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n398_), .B1(new_n419_), .B2(new_n268_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G29gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G43gat), .B(G50gat), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n422_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT15), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G22gat), .ZN(new_n427_));
  INV_X1    g226(.A(G1gat), .ZN(new_n428_));
  INV_X1    g227(.A(G8gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G1gat), .B(G8gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n426_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT76), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n425_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n437_), .A2(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G229gat), .A2(G233gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n437_), .B(new_n433_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT77), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G113gat), .B(G141gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G169gat), .B(G197gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  NOR2_X1   g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n440_), .A2(KEYINPUT77), .A3(new_n443_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n440_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT78), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n450_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G120gat), .B(G148gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT5), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G176gat), .B(G204gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n464_));
  XOR2_X1   g263(.A(G71gat), .B(G78gat), .Z(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n464_), .A2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT12), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n472_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n472_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT7), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n482_), .A2(new_n483_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n472_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n471_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n481_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n487_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT8), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT9), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(G92gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n485_), .A2(KEYINPUT65), .ZN(new_n501_));
  OAI21_X1  g300(.A(G85gat), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n502_), .B2(new_n497_), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT64), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n504_), .A2(new_n507_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n492_), .A2(new_n510_), .A3(new_n489_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT67), .B1(new_n503_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n487_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT9), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n485_), .A2(KEYINPUT65), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n499_), .A2(G92gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n484_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n515_), .B1(new_n518_), .B2(KEYINPUT9), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n479_), .A2(new_n519_), .A3(new_n520_), .A4(new_n510_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n512_), .A2(new_n521_), .A3(KEYINPUT68), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT68), .B1(new_n512_), .B2(new_n521_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n496_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT69), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n496_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n470_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G230gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n512_), .A2(new_n521_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n468_), .B1(new_n496_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n496_), .A2(new_n532_), .A3(new_n468_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(KEYINPUT12), .B2(new_n534_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n528_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n533_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n529_), .B1(new_n537_), .B2(new_n534_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n461_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n536_), .A2(new_n538_), .A3(new_n461_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n457_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT13), .A3(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n420_), .A2(new_n456_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n531_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n512_), .A2(new_n521_), .A3(KEYINPUT68), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n526_), .B1(new_n559_), .B2(new_n496_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n527_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT70), .B(new_n426_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n496_), .A2(new_n532_), .ZN(new_n563_));
  OAI22_X1  g362(.A1(new_n563_), .A2(new_n437_), .B1(KEYINPUT35), .B2(new_n552_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n426_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT70), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n555_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n568_), .A2(KEYINPUT70), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n564_), .B1(new_n568_), .B2(KEYINPUT70), .ZN(new_n572_));
  INV_X1    g371(.A(new_n555_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT71), .ZN(new_n576_));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n570_), .A2(new_n574_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n578_), .B(KEYINPUT36), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n549_), .B(new_n550_), .C1(new_n582_), .C2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n570_), .A2(new_n574_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n583_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n570_), .A2(new_n574_), .A3(new_n581_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n548_), .A3(KEYINPUT37), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n433_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n468_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n594_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT74), .ZN(new_n602_));
  INV_X1    g401(.A(new_n594_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT75), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT75), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n600_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(KEYINPUT74), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n591_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n547_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n356_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n428_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT101), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n588_), .A2(new_n589_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n420_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n609_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n456_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n545_), .A2(new_n620_), .A3(KEYINPUT102), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT102), .B1(new_n545_), .B2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n618_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n428_), .B1(new_n624_), .B2(new_n612_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n614_), .B2(new_n613_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n616_), .A2(new_n626_), .ZN(G1324gat));
  INV_X1    g426(.A(new_n397_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n429_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n624_), .A2(new_n628_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(G8gat), .ZN(new_n632_));
  AOI211_X1 g431(.A(KEYINPUT39), .B(new_n429_), .C1(new_n624_), .C2(new_n628_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g434(.A1(new_n611_), .A2(new_n242_), .A3(new_n268_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n268_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n637_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT41), .B1(new_n637_), .B2(G15gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n638_), .B2(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n611_), .A2(new_n641_), .A3(new_n327_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n624_), .A2(new_n327_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G22gat), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(KEYINPUT42), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(KEYINPUT42), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n617_), .A2(new_n619_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT105), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n547_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(G29gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n612_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n586_), .A2(new_n590_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT103), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n591_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n420_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n658_), .A2(KEYINPUT43), .B1(new_n420_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n623_), .A2(new_n609_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n653_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n661_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n655_), .A2(new_n657_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(new_n420_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n420_), .A2(new_n659_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT44), .B(new_n663_), .C1(new_n666_), .C2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n612_), .A3(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(KEYINPUT104), .ZN(new_n671_));
  OAI21_X1  g470(.A(G29gat), .B1(new_n670_), .B2(KEYINPUT104), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n652_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT106), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n675_), .B(new_n652_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n650_), .A2(new_n678_), .A3(new_n628_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n662_), .A2(new_n628_), .A3(new_n669_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1329gat));
  NAND3_X1  g485(.A1(new_n662_), .A2(new_n268_), .A3(new_n669_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G43gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n650_), .A2(new_n239_), .A3(new_n268_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g490(.A(G50gat), .B1(new_n650_), .B2(new_n327_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n662_), .A2(new_n669_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n327_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(G1331gat));
  NOR3_X1   g494(.A1(new_n546_), .A2(new_n609_), .A3(new_n456_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n618_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n356_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n546_), .A2(new_n456_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n420_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n610_), .ZN(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n612_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n699_), .A2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n706_), .A3(new_n628_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G64gat), .B1(new_n698_), .B2(new_n397_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT48), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT48), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT108), .B(new_n707_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n697_), .B2(new_n268_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT49), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n702_), .A2(new_n716_), .A3(new_n268_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n697_), .B2(new_n327_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT50), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n702_), .A2(new_n721_), .A3(new_n327_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1335gat));
  NAND2_X1  g524(.A1(new_n658_), .A2(KEYINPUT43), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n667_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n700_), .A2(new_n609_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(KEYINPUT109), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n660_), .B2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n356_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n701_), .A2(new_n649_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n484_), .A3(new_n612_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  AOI21_X1  g537(.A(G92gat), .B1(new_n736_), .B2(new_n628_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n397_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n733_), .B2(new_n740_), .ZN(G1337gat));
  INV_X1    g540(.A(G99gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n733_), .B2(new_n268_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n736_), .A2(new_n504_), .A3(new_n508_), .A4(new_n268_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT110), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n744_), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n748_));
  OR2_X1    g547(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n745_), .B(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n748_), .B(new_n749_), .C1(new_n751_), .C2(new_n743_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n747_), .A2(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n727_), .A2(new_n327_), .A3(new_n729_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n759_));
  NOR3_X1   g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n736_), .A2(new_n507_), .A3(new_n509_), .A4(new_n327_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT53), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n758_), .A2(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n756_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n761_), .A4(new_n762_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(G1339gat));
  NAND2_X1  g568(.A1(new_n456_), .A2(new_n543_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n470_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n535_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n529_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n530_), .B1(new_n528_), .B2(new_n535_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(KEYINPUT55), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n772_), .A2(new_n773_), .A3(new_n778_), .A4(new_n529_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n776_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n461_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT56), .B(new_n461_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n770_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n451_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT78), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n436_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n447_), .B1(new_n441_), .B2(new_n439_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n788_), .A2(new_n453_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n543_), .A2(new_n539_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n617_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n543_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n654_), .B1(new_n798_), .B2(KEYINPUT58), .ZN(new_n799_));
  INV_X1    g598(.A(new_n797_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n776_), .A2(new_n779_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT114), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n776_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n461_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n785_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n800_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n799_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT57), .B(new_n617_), .C1(new_n786_), .C2(new_n793_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n796_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n609_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n654_), .A2(new_n619_), .A3(new_n620_), .A4(new_n546_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n268_), .A2(new_n328_), .A3(new_n612_), .A4(new_n397_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT115), .Z(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n456_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n821_), .B(KEYINPUT59), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT116), .B(G113gat), .Z(new_n826_));
  NAND2_X1  g625(.A1(new_n456_), .A2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT117), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n825_), .B2(new_n828_), .ZN(G1340gat));
  XOR2_X1   g628(.A(KEYINPUT118), .B(G120gat), .Z(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n822_), .B(new_n831_), .C1(KEYINPUT60), .C2(new_n830_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n824_), .A2(new_n546_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n830_), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n822_), .B2(new_n619_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n609_), .A2(KEYINPUT119), .ZN(new_n836_));
  MUX2_X1   g635(.A(KEYINPUT119), .B(new_n836_), .S(G127gat), .Z(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n825_), .B2(new_n837_), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n824_), .B2(new_n654_), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n821_), .A2(G134gat), .A3(new_n617_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1343gat));
  NOR4_X1   g640(.A1(new_n268_), .A2(new_n628_), .A3(new_n328_), .A4(new_n356_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n818_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n456_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n546_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT120), .B(G148gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1345gat));
  OR3_X1    g648(.A1(new_n843_), .A2(KEYINPUT121), .A3(new_n609_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT121), .B1(new_n843_), .B2(new_n609_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(new_n617_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G162gat), .B1(new_n844_), .B2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n665_), .A2(G162gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n844_), .B2(new_n858_), .ZN(G1347gat));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n268_), .A2(new_n628_), .A3(new_n356_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n327_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n795_), .A2(new_n794_), .B1(new_n799_), .B2(new_n809_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n619_), .B1(new_n863_), .B2(new_n811_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n456_), .B(new_n862_), .C1(new_n864_), .C2(new_n816_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT62), .B(new_n202_), .C1(new_n865_), .C2(KEYINPUT22), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n816_), .B1(new_n812_), .B2(new_n609_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n862_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n868_), .A2(new_n620_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT22), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G169gat), .B1(new_n865_), .B2(KEYINPUT62), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n860_), .B(new_n866_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n818_), .A2(new_n867_), .A3(new_n456_), .A4(new_n862_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n868_), .A2(KEYINPUT22), .A3(new_n620_), .A4(new_n869_), .ZN(new_n877_));
  OAI211_X1 g676(.A(G169gat), .B(new_n876_), .C1(new_n877_), .C2(new_n867_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n860_), .B1(new_n878_), .B2(new_n866_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n879_), .ZN(G1348gat));
  NOR2_X1   g679(.A1(new_n868_), .A2(new_n869_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G176gat), .B1(new_n881_), .B2(new_n545_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT123), .B1(new_n818_), .B2(new_n328_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n868_), .A2(new_n884_), .A3(new_n327_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n885_), .A3(new_n861_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n546_), .A2(new_n203_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n882_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  AOI21_X1  g687(.A(G183gat), .B1(new_n886_), .B2(new_n619_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n881_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(new_n609_), .A3(new_n213_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n890_), .B2(new_n654_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n617_), .A2(new_n363_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n890_), .B2(new_n894_), .ZN(G1351gat));
  XNOR2_X1  g694(.A(KEYINPUT124), .B(G197gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(G197gat), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n268_), .A2(new_n328_), .A3(new_n612_), .A4(new_n397_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n818_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n620_), .ZN(new_n901_));
  MUX2_X1   g700(.A(new_n896_), .B(new_n898_), .S(new_n901_), .Z(G1352gat));
  AND2_X1   g701(.A1(new_n818_), .A2(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n545_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n619_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n909_));
  INV_X1    g708(.A(G211gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n906_), .A2(KEYINPUT125), .A3(new_n909_), .A4(new_n910_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n908_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  NOR2_X1   g714(.A1(new_n900_), .A2(new_n617_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n916_), .A2(KEYINPUT126), .ZN(new_n917_));
  AOI21_X1  g716(.A(G218gat), .B1(new_n916_), .B2(KEYINPUT126), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n591_), .A2(G218gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT127), .Z(new_n920_));
  AOI22_X1  g719(.A1(new_n917_), .A2(new_n918_), .B1(new_n903_), .B2(new_n920_), .ZN(G1355gat));
endmodule


