//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(KEYINPUT11), .B2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT65), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n202_), .B(new_n206_), .C1(KEYINPUT11), .C2(new_n203_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT66), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT7), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n217_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n224_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT10), .B(G99gat), .Z(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  INV_X1    g033(.A(G92gat), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT9), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n216_), .A2(new_n219_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n229_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n212_), .A2(KEYINPUT12), .A3(new_n240_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G230gat), .A2(G233gat), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n225_), .A2(new_n228_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n211_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n245_), .B2(new_n211_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n244_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n246_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n245_), .A2(new_n211_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n254_));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G176gat), .B(G204gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n249_), .A2(new_n253_), .A3(KEYINPUT68), .A4(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n249_), .A2(new_n253_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n258_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n263_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n263_), .A2(new_n266_), .B1(new_n269_), .B2(new_n267_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT81), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273_));
  INV_X1    g072(.A(G1gat), .ZN(new_n274_));
  INV_X1    g073(.A(G8gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT14), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G8gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G29gat), .B(G36gat), .Z(new_n282_));
  XOR2_X1   g081(.A(G43gat), .B(G50gat), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G29gat), .B(G36gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n287_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n279_), .A2(new_n290_), .A3(new_n280_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(KEYINPUT77), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n281_), .A2(new_n293_), .A3(new_n288_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(G229gat), .A3(G233gat), .A4(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G169gat), .B(G197gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT79), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G141gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n281_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n288_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n290_), .A2(KEYINPUT70), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT15), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(KEYINPUT15), .A3(new_n303_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G229gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT78), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n291_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n295_), .B(new_n299_), .C1(new_n308_), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT80), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n302_), .A2(KEYINPUT15), .A3(new_n303_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT15), .B1(new_n302_), .B2(new_n303_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n281_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n291_), .A3(new_n311_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n295_), .A4(new_n299_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n299_), .B1(new_n318_), .B2(new_n295_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n272_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n272_), .A3(new_n323_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n271_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT85), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT84), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n331_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G71gat), .B(G99gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G183gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT25), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G183gat), .ZN(new_n341_));
  INV_X1    g140(.A(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT26), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G190gat), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n339_), .A2(new_n341_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(G169gat), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(KEYINPUT24), .A3(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n338_), .A2(new_n342_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(KEYINPUT22), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G169gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n366_), .A3(new_n352_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n367_), .A3(new_n354_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n356_), .A2(new_n357_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n357_), .B1(new_n356_), .B2(new_n368_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n356_), .A2(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT82), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n356_), .A2(new_n357_), .A3(new_n368_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT83), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n373_), .A2(new_n378_), .A3(KEYINPUT30), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT30), .B1(new_n373_), .B2(new_n378_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT86), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n371_), .A2(new_n372_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n377_), .A2(KEYINPUT83), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n373_), .A2(new_n378_), .A3(KEYINPUT30), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n337_), .B1(new_n381_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT86), .B1(new_n379_), .B2(new_n380_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n336_), .ZN(new_n391_));
  INV_X1    g190(.A(G134gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G127gat), .ZN(new_n393_));
  INV_X1    g192(.A(G127gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G134gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G120gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G113gat), .ZN(new_n398_));
  INV_X1    g197(.A(G113gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G120gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n393_), .A2(new_n395_), .A3(new_n398_), .A4(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT31), .Z(new_n405_));
  NAND3_X1  g204(.A1(new_n389_), .A2(new_n391_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n386_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n336_), .B1(new_n390_), .B2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n388_), .A2(new_n337_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G155gat), .B(G162gat), .ZN(new_n413_));
  INV_X1    g212(.A(G141gat), .ZN(new_n414_));
  INV_X1    g213(.A(G148gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT3), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(G141gat), .B2(G148gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n413_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(KEYINPUT1), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(new_n415_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G141gat), .A2(G148gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n403_), .B(new_n402_), .C1(new_n423_), .C2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n413_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n416_), .A2(new_n418_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n421_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n433_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n427_), .A2(new_n428_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n429_), .C1(KEYINPUT1), .C2(new_n413_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n440_), .A3(new_n404_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n432_), .A2(new_n441_), .A3(KEYINPUT4), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n432_), .A2(new_n441_), .A3(KEYINPUT97), .A4(KEYINPUT4), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n432_), .B2(KEYINPUT4), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n432_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G1gat), .B(G29gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT0), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G57gat), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n453_), .A2(KEYINPUT0), .ZN(new_n456_));
  INV_X1    g255(.A(G57gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(KEYINPUT0), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n455_), .A2(G85gat), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(G85gat), .B1(new_n455_), .B2(new_n459_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n451_), .A2(new_n452_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n449_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n452_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n438_), .A2(new_n440_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G22gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n472_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G78gat), .B(G106gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT93), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n471_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G211gat), .B(G218gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482_));
  INV_X1    g281(.A(G204gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(G197gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(G197gat), .ZN(new_n485_));
  INV_X1    g284(.A(G197gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n488_), .B2(KEYINPUT21), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT88), .B1(new_n483_), .B2(G197gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n486_), .A3(G204gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n492_), .A3(new_n485_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT21), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT89), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n496_), .A3(KEYINPUT21), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n489_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n481_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT21), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n488_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n484_), .A2(new_n487_), .A3(KEYINPUT91), .A4(new_n485_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n480_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT92), .B1(new_n498_), .B2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G228gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n499_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n493_), .A2(new_n496_), .A3(KEYINPUT21), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n496_), .B1(new_n493_), .B2(KEYINPUT21), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n502_), .A2(new_n503_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(KEYINPUT21), .A3(new_n499_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n479_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n520_), .B2(new_n507_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n478_), .B1(new_n509_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n476_), .B1(new_n522_), .B2(KEYINPUT94), .ZN(new_n523_));
  INV_X1    g322(.A(new_n478_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n518_), .A2(new_n520_), .A3(new_n507_), .ZN(new_n525_));
  AOI221_X4 g324(.A(new_n479_), .B1(new_n519_), .B2(new_n508_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n509_), .A2(new_n521_), .A3(new_n478_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n527_), .A2(KEYINPUT94), .A3(new_n528_), .A4(new_n476_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n515_), .A2(new_n517_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n377_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT19), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n356_), .A2(new_n368_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n515_), .A2(new_n517_), .A3(new_n540_), .A4(KEYINPUT95), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n515_), .A2(new_n517_), .A3(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n536_), .A2(new_n539_), .A3(new_n541_), .A4(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n375_), .A2(new_n515_), .A3(new_n517_), .A4(new_n376_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n374_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(KEYINPUT20), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n538_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G8gat), .B(G36gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n545_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n533_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n539_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n546_), .A2(new_n547_), .A3(KEYINPUT20), .A4(new_n539_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n554_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n545_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(KEYINPUT27), .A3(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n558_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n412_), .A2(new_n470_), .A3(new_n532_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n530_), .A2(new_n531_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n470_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n495_), .A2(new_n497_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n504_), .B1(new_n570_), .B2(new_n512_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT20), .B(new_n542_), .C1(new_n371_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n538_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n560_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n555_), .A2(KEYINPUT32), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n545_), .A2(new_n549_), .A3(new_n575_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n468_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n464_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n466_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT33), .A3(new_n463_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n461_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n455_), .A2(G85gat), .A3(new_n459_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n432_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n432_), .A2(KEYINPUT4), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n448_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n446_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(new_n583_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n545_), .A2(new_n549_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n554_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n563_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n579_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n532_), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n567_), .B(new_n412_), .C1(new_n569_), .C2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT33), .B1(new_n582_), .B2(new_n463_), .ZN(new_n599_));
  NOR4_X1   g398(.A1(new_n465_), .A2(new_n580_), .A3(new_n466_), .A4(new_n462_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n590_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n556_), .A2(new_n557_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n467_), .A2(new_n464_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n601_), .A2(new_n602_), .B1(new_n603_), .B2(new_n578_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n558_), .A2(new_n531_), .A3(new_n530_), .A4(new_n564_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n468_), .A2(new_n469_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT98), .B1(new_n464_), .B2(new_n467_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n604_), .A2(new_n568_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n406_), .A2(new_n411_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT100), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n566_), .B1(new_n598_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(G183gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT76), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n212_), .A2(new_n242_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT74), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n281_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n620_), .B(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n616_), .B(KEYINPUT17), .Z(new_n626_));
  XOR2_X1   g425(.A(new_n623_), .B(new_n211_), .Z(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n240_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT34), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n245_), .A2(new_n290_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n631_), .B(new_n636_), .C1(new_n632_), .C2(new_n635_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G190gat), .B(G218gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(KEYINPUT36), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n639_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT71), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n640_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n643_), .B(KEYINPUT36), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT72), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n649_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT73), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(KEYINPUT37), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(KEYINPUT37), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n647_), .A2(new_n648_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n656_), .A3(KEYINPUT37), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  AND4_X1   g462(.A1(new_n329_), .A2(new_n612_), .A3(new_n630_), .A4(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n274_), .A3(new_n608_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n661_), .B(new_n668_), .ZN(new_n669_));
  AND4_X1   g468(.A1(new_n329_), .A2(new_n612_), .A3(new_n630_), .A4(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n274_), .B1(new_n670_), .B2(new_n608_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n667_), .A2(new_n671_), .ZN(G1324gat));
  INV_X1    g471(.A(new_n565_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n275_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n673_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(G8gat), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n675_), .B2(G8gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT104), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n681_), .B(new_n674_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n680_), .A2(KEYINPUT40), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT40), .B1(new_n680_), .B2(new_n682_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n670_), .B2(new_n412_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT41), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n664_), .A2(new_n686_), .A3(new_n412_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1326gat));
  INV_X1    g489(.A(G22gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n670_), .B2(new_n568_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT42), .Z(new_n693_));
  NAND2_X1  g492(.A1(new_n568_), .A2(new_n691_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n664_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n655_), .A2(new_n630_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n612_), .A2(new_n329_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G29gat), .B1(new_n699_), .B2(new_n608_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n329_), .A2(new_n629_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n566_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n605_), .A2(new_n608_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n590_), .B1(new_n464_), .B2(new_n580_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(new_n563_), .A3(new_n594_), .A4(new_n583_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n705_), .A2(new_n579_), .B1(new_n531_), .B2(new_n530_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n610_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n567_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n609_), .A2(KEYINPUT100), .A3(new_n610_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n702_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n710_), .B2(new_n663_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n660_), .A2(new_n662_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n612_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n701_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT44), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n716_), .A2(G29gat), .A3(new_n608_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n701_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n710_), .A2(KEYINPUT43), .A3(new_n663_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n712_), .B1(new_n612_), .B2(new_n713_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n700_), .B1(new_n717_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n699_), .A2(new_n725_), .A3(new_n673_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n565_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n723_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(G36gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT106), .B(new_n725_), .C1(new_n729_), .C2(new_n723_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT46), .B(new_n727_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  NAND3_X1  g536(.A1(new_n716_), .A2(G43gat), .A3(new_n412_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n723_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n699_), .A2(new_n412_), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n738_), .A2(new_n739_), .B1(G43gat), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n699_), .B2(new_n568_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n716_), .A2(G50gat), .A3(new_n568_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n723_), .ZN(G1331gat));
  AND3_X1   g544(.A1(new_n612_), .A2(KEYINPUT107), .A3(new_n328_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT107), .B1(new_n612_), .B2(new_n328_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n271_), .ZN(new_n749_));
  NOR4_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n629_), .A4(new_n713_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT108), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n457_), .A3(new_n608_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n669_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n710_), .A2(new_n753_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n749_), .A2(new_n327_), .A3(new_n629_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n470_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n752_), .A2(new_n758_), .ZN(G1332gat));
  INV_X1    g558(.A(G64gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n751_), .A2(new_n760_), .A3(new_n673_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G64gat), .B1(new_n757_), .B2(new_n565_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT109), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT109), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(KEYINPUT48), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT48), .B1(new_n763_), .B2(new_n764_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n751_), .A2(new_n768_), .A3(new_n412_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n756_), .B2(new_n412_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT49), .Z(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1334gat));
  INV_X1    g571(.A(G78gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n751_), .A2(new_n773_), .A3(new_n568_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n756_), .B2(new_n568_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT50), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1335gat));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n711_), .A2(new_n714_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n749_), .A2(new_n327_), .A3(new_n630_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n780_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n778_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT111), .A3(new_n782_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(G85gat), .A4(new_n608_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n271_), .B(new_n698_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n234_), .B1(new_n790_), .B2(new_n470_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT112), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(new_n794_), .A3(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1336gat));
  NAND4_X1  g595(.A1(new_n785_), .A2(new_n788_), .A3(G92gat), .A4(new_n673_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n235_), .B1(new_n790_), .B2(new_n565_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1337gat));
  INV_X1    g598(.A(new_n790_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n230_), .A3(new_n412_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n610_), .B1(new_n787_), .B2(new_n782_), .ZN(new_n802_));
  INV_X1    g601(.A(G99gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g604(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n790_), .A2(G106gat), .A3(new_n532_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G106gat), .B1(new_n786_), .B2(new_n532_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT52), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT52), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n807_), .B(new_n808_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n809_), .B(KEYINPUT52), .ZN(new_n813_));
  INV_X1    g612(.A(new_n808_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n806_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n812_), .A2(new_n815_), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n263_), .A2(new_n266_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n317_), .A2(new_n291_), .A3(new_n310_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n299_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n292_), .A2(new_n294_), .A3(new_n311_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n321_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n823_), .A2(new_n828_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT81), .B(new_n322_), .C1(new_n314_), .C2(new_n320_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n263_), .B1(new_n830_), .B2(new_n324_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n249_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n249_), .A2(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n249_), .A2(KEYINPUT115), .A3(new_n832_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n243_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n250_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .A4(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n840_), .B2(new_n265_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n831_), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n832_), .B2(new_n249_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT115), .B1(new_n249_), .B2(new_n832_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n258_), .B1(new_n846_), .B2(new_n837_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n847_), .B2(KEYINPUT116), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n829_), .B1(new_n842_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n661_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n822_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n829_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n249_), .A2(KEYINPUT115), .A3(new_n832_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n844_), .A2(new_n855_), .A3(new_n845_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n854_), .B(KEYINPUT56), .C1(new_n856_), .C2(new_n258_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n325_), .A2(new_n326_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n841_), .A2(KEYINPUT56), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n853_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n821_), .A3(new_n850_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n843_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n863_), .B(new_n865_), .C1(new_n856_), .C2(new_n258_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n840_), .A2(new_n864_), .A3(new_n843_), .A4(new_n265_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n828_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n866_), .A2(KEYINPUT58), .A3(new_n867_), .A4(new_n868_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n713_), .A3(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n852_), .A2(new_n862_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n629_), .ZN(new_n875_));
  AND2_X1   g674(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n327_), .A2(new_n629_), .A3(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n663_), .A2(new_n749_), .A3(new_n877_), .A4(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n877_), .B1(new_n270_), .B2(new_n268_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n881_), .B2(new_n713_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n568_), .B1(new_n875_), .B2(new_n884_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n610_), .A2(new_n673_), .A3(new_n470_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n818_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n874_), .B2(new_n629_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n886_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n888_), .A2(KEYINPUT59), .A3(new_n568_), .A4(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n327_), .A2(G113gat), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n887_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n888_), .A2(new_n568_), .A3(new_n889_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G113gat), .B1(new_n893_), .B2(new_n327_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n817_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n875_), .A2(new_n884_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n532_), .A3(new_n886_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n399_), .B1(new_n897_), .B2(new_n328_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(KEYINPUT59), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n885_), .A2(new_n818_), .A3(new_n886_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT119), .B(new_n898_), .C1(new_n901_), .C2(new_n891_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n895_), .A2(new_n902_), .ZN(G1340gat));
  OAI21_X1  g702(.A(G120gat), .B1(new_n901_), .B2(new_n749_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905_));
  AOI21_X1  g704(.A(G120gat), .B1(new_n271_), .B2(new_n905_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT120), .Z(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n905_), .B2(G120gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n893_), .A2(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT121), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n904_), .A2(new_n910_), .ZN(G1341gat));
  NAND2_X1  g710(.A1(new_n630_), .A2(G127gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n887_), .A2(new_n890_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G127gat), .B1(new_n893_), .B2(new_n630_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n394_), .B1(new_n897_), .B2(new_n629_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n916_), .B(new_n917_), .C1(new_n901_), .C2(new_n912_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n918_), .ZN(G1342gat));
  INV_X1    g718(.A(new_n901_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n663_), .A2(new_n392_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n392_), .B1(new_n897_), .B2(new_n669_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT123), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n924_), .B(new_n392_), .C1(new_n897_), .C2(new_n669_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n920_), .A2(new_n921_), .B1(new_n923_), .B2(new_n925_), .ZN(G1343gat));
  NOR3_X1   g725(.A1(new_n412_), .A2(new_n470_), .A3(new_n605_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n896_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n328_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n414_), .ZN(G1344gat));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n749_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n415_), .ZN(G1345gat));
  NOR2_X1   g731(.A1(new_n928_), .A2(new_n629_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT61), .B(G155gat), .Z(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1346gat));
  INV_X1    g734(.A(G162gat), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n928_), .A2(new_n936_), .A3(new_n663_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n928_), .B2(new_n669_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n939_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n937_), .B1(new_n940_), .B2(new_n941_), .ZN(G1347gat));
  INV_X1    g741(.A(new_n885_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n412_), .A2(new_n470_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n565_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n943_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n327_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n943_), .A2(new_n328_), .A3(new_n946_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n950_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n950_), .B2(new_n351_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n949_), .A2(new_n951_), .A3(new_n953_), .ZN(G1348gat));
  NAND2_X1  g753(.A1(new_n947_), .A2(new_n271_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g755(.A(G183gat), .B1(new_n947_), .B2(new_n630_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n339_), .A2(new_n341_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n885_), .A2(new_n630_), .A3(new_n958_), .A4(new_n945_), .ZN(new_n959_));
  AND2_X1   g758(.A1(new_n959_), .A2(KEYINPUT125), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n959_), .A2(KEYINPUT125), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n957_), .A2(new_n960_), .A3(new_n961_), .ZN(G1350gat));
  NAND4_X1  g761(.A1(new_n947_), .A2(new_n753_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n943_), .A2(new_n663_), .A3(new_n946_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n342_), .ZN(G1351gat));
  NOR3_X1   g764(.A1(new_n412_), .A2(new_n608_), .A3(new_n532_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n966_), .A2(new_n967_), .ZN(new_n969_));
  NOR4_X1   g768(.A1(new_n888_), .A2(new_n565_), .A3(new_n968_), .A4(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n327_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n271_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g773(.A1(new_n970_), .A2(new_n630_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  AND2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n975_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n978_), .B1(new_n975_), .B2(new_n976_), .ZN(G1354gat));
  INV_X1    g778(.A(G218gat), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n970_), .A2(new_n980_), .A3(new_n753_), .ZN(new_n981_));
  AND2_X1   g780(.A1(new_n970_), .A2(new_n713_), .ZN(new_n982_));
  OAI211_X1 g781(.A(KEYINPUT127), .B(new_n981_), .C1(new_n982_), .C2(new_n980_), .ZN(new_n983_));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984_));
  AND3_X1   g783(.A1(new_n970_), .A2(new_n980_), .A3(new_n753_), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n980_), .B1(new_n970_), .B2(new_n713_), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n984_), .B1(new_n985_), .B2(new_n986_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n983_), .A2(new_n987_), .ZN(G1355gat));
endmodule


