//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT8), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT7), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n205_), .A2(new_n214_), .A3(new_n206_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n208_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G92gat), .Z(new_n217_));
  NOR3_X1   g016(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n203_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n205_), .A2(new_n219_), .ZN(new_n220_));
  OAI22_X1  g019(.A1(new_n218_), .A2(new_n220_), .B1(G85gat), .B2(G92gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n221_), .A2(new_n224_), .B1(new_n214_), .B2(new_n210_), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n212_), .B(KEYINPUT65), .Z(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT66), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(new_n232_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n235_), .B(KEYINPUT68), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n228_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n227_), .A2(KEYINPUT12), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n227_), .B(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT12), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G230gat), .A2(G233gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n247_), .A2(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n244_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(G230gat), .A3(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G120gat), .B(G148gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT5), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT69), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n256_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT70), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n253_), .A2(new_n256_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(new_n262_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT13), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n266_), .A2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n202_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n266_), .A2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n267_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT71), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G1gat), .ZN(new_n275_));
  INV_X1    g074(.A(G8gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT74), .B(G15gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n279_), .B2(G22gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(G22gat), .B2(new_n279_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G1gat), .B(G8gat), .Z(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G43gat), .B(G50gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n283_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G229gat), .A2(G233gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n286_), .B(KEYINPUT15), .ZN(new_n290_));
  MUX2_X1   g089(.A(new_n290_), .B(new_n286_), .S(new_n283_), .Z(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G113gat), .B(G141gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G169gat), .B(G197gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n292_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n274_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G71gat), .B(G99gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT78), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G227gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G43gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT77), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n303_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT23), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  INV_X1    g111(.A(G176gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT26), .B(G190gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT25), .B(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT26), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n317_), .B1(new_n320_), .B2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n308_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n313_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n325_), .A2(KEYINPUT24), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT24), .A3(new_n310_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n315_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT30), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n306_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT31), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333_));
  XOR2_X1   g132(.A(G113gat), .B(G120gat), .Z(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n335_), .A2(KEYINPUT79), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(KEYINPUT79), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n334_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n332_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n307_), .B(KEYINPUT23), .Z(new_n351_));
  INV_X1    g150(.A(new_n322_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT26), .B(G190gat), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT76), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n328_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n355_), .A2(new_n356_), .B1(new_n314_), .B2(new_n309_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(G211gat), .B(G218gat), .Z(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT21), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT86), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n358_), .A3(KEYINPUT21), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n357_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT20), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n366_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n314_), .A2(KEYINPUT92), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n314_), .A2(KEYINPUT92), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n309_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n316_), .A2(new_n319_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n356_), .A2(new_n308_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n370_), .A2(KEYINPUT91), .B1(new_n371_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(new_n379_), .A3(KEYINPUT20), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n350_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n371_), .A2(KEYINPUT86), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n329_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n371_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n376_), .A3(new_n374_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n349_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n347_), .B1(new_n381_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n329_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT91), .B1(new_n392_), .B2(new_n387_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n377_), .A2(new_n371_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n380_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n390_), .B1(new_n395_), .B2(new_n349_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n346_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n400_));
  NAND3_X1  g199(.A1(new_n384_), .A2(new_n386_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n349_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n395_), .B2(new_n349_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n346_), .B(KEYINPUT97), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n399_), .B1(new_n396_), .B2(new_n346_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n398_), .A2(new_n399_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n342_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT80), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(G141gat), .A3(G148gat), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G141gat), .A2(G148gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT81), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(KEYINPUT1), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n420_), .B2(KEYINPUT1), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(KEYINPUT83), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n428_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR4_X1   g229(.A1(KEYINPUT82), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n416_), .B2(new_n433_), .ZN(new_n434_));
  OAI22_X1  g233(.A1(new_n427_), .A2(new_n430_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT2), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n412_), .A2(new_n414_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n425_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n437_), .A2(new_n438_), .ZN(new_n441_));
  INV_X1    g240(.A(G141gat), .ZN(new_n442_));
  INV_X1    g241(.A(G148gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n433_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT82), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n416_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n426_), .A2(KEYINPUT83), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n445_), .A2(new_n446_), .B1(new_n447_), .B2(new_n429_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n441_), .A2(new_n448_), .A3(KEYINPUT84), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n420_), .B1(G155gat), .B2(G162gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n424_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT29), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n382_), .A2(new_n383_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT85), .Z(new_n458_));
  NOR3_X1   g257(.A1(new_n455_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT87), .B1(new_n453_), .B2(new_n454_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n451_), .B1(new_n440_), .B2(new_n449_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n461_), .B(KEYINPUT29), .C1(new_n462_), .C2(new_n424_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n464_), .B2(new_n371_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n465_), .B2(KEYINPUT88), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n385_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n457_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n410_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n435_), .A2(new_n425_), .A3(new_n439_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT84), .B1(new_n441_), .B2(new_n448_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n452_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n424_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n461_), .B1(new_n475_), .B2(KEYINPUT29), .ZN(new_n476_));
  INV_X1    g275(.A(new_n463_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n371_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n457_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(KEYINPUT88), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n459_), .ZN(new_n481_));
  AND4_X1   g280(.A1(new_n469_), .A2(new_n480_), .A3(new_n481_), .A4(new_n410_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT90), .B1(new_n470_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n453_), .A2(new_n454_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G22gat), .B(G50gat), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n486_), .B(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n480_), .A2(new_n469_), .A3(new_n481_), .A4(new_n410_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n480_), .A2(new_n469_), .A3(new_n481_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n409_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n490_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n483_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n483_), .B2(new_n496_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n475_), .A2(new_n340_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n473_), .B(new_n474_), .C1(new_n335_), .C2(new_n339_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n501_), .A2(KEYINPUT4), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n501_), .B2(KEYINPUT4), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n502_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n503_), .A2(new_n506_), .B1(new_n507_), .B2(new_n505_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G29gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT0), .ZN(new_n511_));
  INV_X1    g310(.A(G57gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(new_n203_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n508_), .A2(new_n509_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  OAI221_X1 g315(.A(new_n516_), .B1(new_n507_), .B2(new_n505_), .C1(new_n503_), .C2(new_n506_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n509_), .B1(new_n508_), .B2(new_n514_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n500_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n508_), .A2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT95), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(KEYINPUT96), .A3(new_n515_), .A4(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n408_), .A2(new_n499_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n407_), .A3(new_n523_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n497_), .A2(new_n498_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n501_), .A2(KEYINPUT4), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT4), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n504_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT93), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n528_), .A2(new_n532_), .A3(new_n504_), .A4(new_n529_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n507_), .A2(new_n504_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n516_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n531_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(new_n398_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n517_), .B(KEYINPUT33), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n522_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n381_), .A2(new_n540_), .A3(new_n390_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n403_), .B2(new_n540_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n537_), .A2(new_n538_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n492_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n470_), .A2(new_n482_), .A3(KEYINPUT90), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n495_), .B1(new_n494_), .B2(new_n490_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n483_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n341_), .B1(new_n527_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT98), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n537_), .A2(new_n538_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n539_), .A2(new_n542_), .ZN(new_n553_));
  OAI22_X1  g352(.A1(new_n497_), .A2(new_n498_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n520_), .A2(new_n407_), .A3(new_n523_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n547_), .A2(new_n555_), .A3(new_n548_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n341_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n525_), .B1(new_n551_), .B2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n299_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n228_), .A2(new_n286_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT35), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n227_), .A2(new_n290_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n563_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n570_), .A2(KEYINPUT36), .A3(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(KEYINPUT36), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n578_));
  NOR2_X1   g377(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n283_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n243_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n582_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n561_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n275_), .A3(new_n524_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT38), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n577_), .B(KEYINPUT99), .ZN(new_n600_));
  NOR4_X1   g399(.A1(new_n299_), .A2(new_n560_), .A3(new_n600_), .A4(new_n595_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n524_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(new_n407_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n276_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n606_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(G8gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n608_), .B2(G8gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT100), .B(new_n609_), .C1(new_n608_), .C2(G8gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT40), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT40), .B(new_n607_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1325gat));
  OAI21_X1  g418(.A(G15gat), .B1(new_n602_), .B2(new_n341_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT41), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT41), .ZN(new_n622_));
  INV_X1    g421(.A(G15gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n597_), .A2(new_n623_), .A3(new_n342_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n621_), .A2(new_n622_), .A3(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n601_), .B2(new_n499_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT42), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n597_), .A2(new_n626_), .A3(new_n499_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n595_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n577_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n561_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n524_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n298_), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n636_), .B(new_n631_), .C1(new_n270_), .C2(new_n273_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n582_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT101), .B(KEYINPUT43), .C1(new_n560_), .C2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n525_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n558_), .B1(new_n557_), .B2(new_n341_), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT98), .B(new_n342_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n582_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n582_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT101), .B1(new_n647_), .B2(KEYINPUT43), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n637_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT44), .B(new_n637_), .C1(new_n646_), .C2(new_n648_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n524_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n635_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  NOR2_X1   g454(.A1(new_n407_), .A2(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n561_), .A2(new_n632_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n651_), .A2(new_n606_), .A3(new_n652_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n659_), .A2(KEYINPUT102), .A3(G36gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT102), .B1(new_n659_), .B2(G36gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(KEYINPUT46), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  OAI221_X1 g464(.A(new_n658_), .B1(new_n663_), .B2(KEYINPUT46), .C1(new_n660_), .C2(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1329gat));
  INV_X1    g466(.A(G43gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n341_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n651_), .A2(new_n652_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n651_), .A2(KEYINPUT104), .A3(new_n652_), .A4(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n668_), .B1(new_n633_), .B2(new_n341_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n634_), .B2(new_n499_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n499_), .A2(G50gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n653_), .B2(new_n682_), .ZN(G1331gat));
  INV_X1    g482(.A(new_n274_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n596_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n636_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n686_), .B2(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n643_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(G57gat), .A3(new_n603_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n595_), .A2(new_n298_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n560_), .A3(new_n600_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n512_), .B1(new_n693_), .B2(new_n524_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n606_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(G64gat), .ZN(new_n698_));
  INV_X1    g497(.A(G64gat), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT48), .B(new_n699_), .C1(new_n693_), .C2(new_n606_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n606_), .A2(new_n699_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n698_), .A2(new_n700_), .B1(new_n689_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n693_), .B2(new_n342_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT49), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n342_), .A2(new_n704_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n689_), .B2(new_n707_), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n693_), .A2(new_n499_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G78gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n711_));
  OR2_X1    g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n711_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n497_), .A2(new_n498_), .A3(G78gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT108), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n688_), .A2(new_n643_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n712_), .A2(KEYINPUT109), .A3(new_n713_), .A4(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1335gat));
  NAND2_X1  g520(.A1(new_n684_), .A2(new_n636_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n577_), .A3(new_n631_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n643_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n203_), .B1(new_n724_), .B2(new_n603_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n646_), .A2(new_n648_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n722_), .A2(new_n631_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n524_), .A2(G85gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT110), .Z(new_n730_));
  OAI21_X1  g529(.A(new_n725_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT111), .Z(G1336gat));
  OAI21_X1  g531(.A(new_n204_), .B1(new_n724_), .B2(new_n407_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n407_), .A2(new_n217_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n728_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT112), .ZN(G1337gat));
  OAI21_X1  g535(.A(G99gat), .B1(new_n728_), .B2(new_n341_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n342_), .A2(new_n222_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n724_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n726_), .A2(new_n499_), .A3(new_n727_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G106gat), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n499_), .A2(new_n223_), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n743_), .A2(new_n744_), .B1(new_n724_), .B2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(G1339gat));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n253_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n251_), .A2(KEYINPUT55), .A3(new_n252_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n750_), .B(new_n751_), .C1(new_n252_), .C2(new_n251_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(KEYINPUT56), .A3(new_n261_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT56), .B1(new_n752_), .B2(new_n261_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n754_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n292_), .A2(new_n295_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n291_), .A2(new_n288_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n288_), .B2(new_n287_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n295_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n264_), .A2(new_n765_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n760_), .A2(new_n761_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n761_), .B1(new_n760_), .B2(new_n766_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n582_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n756_), .A2(KEYINPUT115), .A3(new_n753_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n752_), .A2(new_n771_), .A3(KEYINPUT56), .A4(new_n261_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(new_n298_), .A3(new_n264_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT116), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n773_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n266_), .A2(new_n765_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT57), .A3(new_n577_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n769_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT57), .B1(new_n779_), .B2(new_n577_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n595_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n266_), .B(KEYINPUT13), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n691_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n638_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n785_), .B2(new_n691_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n784_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT54), .A3(new_n638_), .A4(new_n787_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n603_), .B1(new_n783_), .B2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n408_), .A2(new_n499_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT118), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n798_), .A3(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(new_n298_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(G113gat), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n794_), .A2(KEYINPUT59), .A3(new_n795_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n298_), .A2(new_n806_), .A3(G113gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n806_), .B2(G113gat), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n800_), .A2(new_n801_), .B1(new_n805_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n810_));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n684_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n797_), .A2(new_n799_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n274_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n811_), .ZN(G1341gat));
  NAND3_X1  g615(.A1(new_n797_), .A2(new_n631_), .A3(new_n799_), .ZN(new_n817_));
  INV_X1    g616(.A(G127gat), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n631_), .A2(new_n819_), .A3(G127gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n819_), .B2(G127gat), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n817_), .A2(new_n818_), .B1(new_n805_), .B2(new_n821_), .ZN(G1342gat));
  NAND3_X1  g621(.A1(new_n797_), .A2(new_n600_), .A3(new_n799_), .ZN(new_n823_));
  INV_X1    g622(.A(G134gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n582_), .A2(G134gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT121), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n823_), .A2(new_n824_), .B1(new_n805_), .B2(new_n826_), .ZN(G1343gat));
  NAND2_X1  g626(.A1(new_n499_), .A2(new_n341_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n606_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n794_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n636_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT122), .B(G141gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n830_), .A2(new_n274_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT123), .B(G148gat), .Z(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1345gat));
  NAND2_X1  g635(.A1(new_n783_), .A2(new_n793_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n837_), .A2(new_n524_), .A3(new_n631_), .A4(new_n829_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n794_), .A2(KEYINPUT124), .A3(new_n631_), .A4(new_n829_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1346gat));
  INV_X1    g644(.A(new_n830_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G162gat), .B1(new_n846_), .B2(new_n600_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n582_), .A2(G162gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT125), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n846_), .B2(new_n849_), .ZN(G1347gat));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n603_), .A2(new_n606_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n499_), .A2(new_n852_), .A3(new_n341_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n837_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n636_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n851_), .B1(new_n855_), .B2(new_n324_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT62), .B(G169gat), .C1(new_n854_), .C2(new_n636_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n312_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(G1348gat));
  NOR2_X1   g658(.A1(new_n854_), .A2(new_n274_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n313_), .ZN(G1349gat));
  NOR2_X1   g660(.A1(new_n854_), .A2(new_n595_), .ZN(new_n862_));
  MUX2_X1   g661(.A(G183gat), .B(new_n319_), .S(new_n862_), .Z(G1350gat));
  OAI21_X1  g662(.A(G190gat), .B1(new_n854_), .B2(new_n638_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n600_), .A2(new_n316_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n854_), .B2(new_n865_), .ZN(G1351gat));
  INV_X1    g665(.A(G197gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n828_), .A2(new_n852_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n837_), .A2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(KEYINPUT126), .B(new_n867_), .C1(new_n869_), .C2(new_n636_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n837_), .A2(new_n868_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n298_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n872_), .B2(new_n867_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n867_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1352gat));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n684_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g676(.A(KEYINPUT63), .B(G211gat), .Z(new_n878_));
  NAND4_X1  g677(.A1(new_n871_), .A2(KEYINPUT127), .A3(new_n631_), .A4(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n869_), .A2(new_n595_), .ZN(new_n880_));
  OR2_X1    g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT127), .B1(new_n880_), .B2(new_n878_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1354gat));
  INV_X1    g683(.A(G218gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n871_), .A2(new_n885_), .A3(new_n600_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G218gat), .B1(new_n869_), .B2(new_n638_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1355gat));
endmodule


