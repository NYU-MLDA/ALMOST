//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n203_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(new_n206_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT12), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n216_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G85gat), .B(G92gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n227_), .A3(new_n224_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT8), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(KEYINPUT64), .ZN(new_n230_));
  AND3_X1   g029(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n221_), .A4(new_n216_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n230_), .A2(new_n235_), .A3(new_n236_), .A4(new_n224_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT9), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(G85gat), .A3(G92gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n233_), .B(new_n240_), .C1(new_n239_), .C2(new_n223_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT10), .B(G99gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(G106gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT67), .B1(new_n238_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  AOI211_X1 g046(.A(new_n247_), .B(new_n244_), .C1(new_n229_), .C2(new_n237_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n212_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n222_), .A2(new_n227_), .A3(new_n224_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n227_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n236_), .ZN(new_n252_));
  AND4_X1   g051(.A1(new_n236_), .A2(new_n230_), .A3(new_n235_), .A4(new_n224_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n245_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n205_), .A2(new_n206_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n202_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n208_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n207_), .B2(new_n209_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n211_), .ZN(new_n262_));
  AND2_X1   g061(.A1(G230gat), .A2(G233gat), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n258_), .A2(new_n259_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n244_), .B1(new_n229_), .B2(new_n237_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n249_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT68), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n249_), .A2(new_n262_), .A3(new_n266_), .A4(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n264_), .A2(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n261_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n263_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n271_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT69), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(KEYINPUT69), .ZN(new_n284_));
  OAI22_X1  g083(.A1(new_n280_), .A2(new_n281_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n281_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n271_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n288_), .B2(new_n283_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G43gat), .B(G50gat), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n298_), .B(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n298_), .A2(new_n305_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT15), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n305_), .B(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n309_), .B2(new_n298_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311_));
  MUX2_X1   g110(.A(new_n306_), .B(new_n310_), .S(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G169gat), .B(G197gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n312_), .B(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n289_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n324_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326_));
  INV_X1    g125(.A(G141gat), .ZN(new_n327_));
  INV_X1    g126(.A(G148gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .A4(KEYINPUT84), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n323_), .A2(KEYINPUT85), .A3(new_n325_), .A4(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n329_), .A2(new_n325_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n330_), .A2(new_n333_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n327_), .A2(new_n328_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n319_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G127gat), .A2(G134gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G127gat), .A2(G134gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(G120gat), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G120gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n343_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT82), .B(G113gat), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n342_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n336_), .A2(new_n353_), .A3(new_n341_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT4), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT96), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n355_), .A2(new_n358_), .A3(KEYINPUT4), .A4(new_n356_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n318_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n356_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(new_n359_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n318_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n364_), .A2(new_n368_), .A3(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT33), .B1(new_n374_), .B2(KEYINPUT97), .ZN(new_n375_));
  XOR2_X1   g174(.A(G64gat), .B(G92gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT23), .ZN(new_n383_));
  OR2_X1    g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(KEYINPUT24), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n388_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n383_), .B1(G183gat), .B2(G190gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT22), .B(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n386_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G197gat), .A2(G204gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT88), .B(G197gat), .Z(new_n402_));
  OAI211_X1 g201(.A(KEYINPUT21), .B(new_n401_), .C1(new_n402_), .C2(G204gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n404_));
  INV_X1    g203(.A(G204gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G197gat), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n404_), .B(new_n406_), .C1(new_n402_), .C2(new_n405_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n406_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n408_), .A2(KEYINPUT90), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(KEYINPUT90), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(KEYINPUT21), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT20), .B1(new_n400_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G183gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(G183gat), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n392_), .B(new_n417_), .C1(new_n418_), .C2(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n388_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n383_), .B1(G190gat), .B2(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n398_), .A2(KEYINPUT81), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n396_), .A2(new_n423_), .A3(new_n397_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n386_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(new_n414_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n415_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n400_), .B2(new_n414_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n420_), .A2(new_n425_), .A3(new_n409_), .A4(new_n413_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n430_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n381_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n415_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n427_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n430_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n400_), .A2(new_n414_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT20), .A3(new_n435_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n431_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n443_), .A3(new_n380_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n318_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n366_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n362_), .A2(new_n363_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n372_), .B1(new_n448_), .B2(new_n318_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n446_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n375_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n431_), .B1(new_n415_), .B2(new_n427_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n434_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n440_), .A2(new_n443_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n372_), .B1(new_n451_), .B2(new_n367_), .ZN(new_n463_));
  OAI221_X1 g262(.A(new_n461_), .B1(new_n460_), .B2(new_n462_), .C1(new_n463_), .C2(new_n374_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n420_), .A2(new_n425_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n426_), .A2(KEYINPUT30), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G43gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G71gat), .B(G99gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n353_), .A2(KEYINPUT31), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n353_), .A2(KEYINPUT31), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n480_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n472_), .A2(new_n474_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n477_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n486_), .B1(new_n490_), .B2(new_n479_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n414_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n409_), .A2(new_n413_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT91), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G233gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(KEYINPUT87), .A2(G228gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT87), .A2(G228gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n497_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n494_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n513_));
  OR3_X1    g312(.A1(new_n342_), .A2(KEYINPUT29), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G22gat), .B(G50gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n342_), .B2(KEYINPUT29), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n515_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n512_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n516_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT92), .A3(new_n517_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n497_), .A2(new_n501_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n506_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n494_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n508_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n511_), .A2(new_n520_), .A3(new_n524_), .A4(new_n528_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n518_), .A2(new_n519_), .A3(new_n512_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n509_), .A2(new_n510_), .A3(new_n494_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n526_), .B2(new_n508_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n493_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n465_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n463_), .A2(new_n374_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n444_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n380_), .B(KEYINPUT98), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT27), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n537_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT27), .B1(new_n437_), .B2(new_n444_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n533_), .A2(new_n492_), .A3(new_n529_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n492_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n536_), .B(new_n543_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n535_), .A2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n317_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G190gat), .B(G218gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  INV_X1    g352(.A(new_n305_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n245_), .B(new_n554_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n265_), .A2(KEYINPUT72), .A3(new_n554_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n309_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT70), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n562_), .B(new_n563_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n557_), .A2(new_n561_), .A3(new_n564_), .A4(new_n560_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n309_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n254_), .A2(new_n247_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n265_), .A2(KEYINPUT67), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n569_), .B(new_n566_), .C1(new_n570_), .C2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n553_), .B1(new_n568_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n552_), .B1(new_n576_), .B2(new_n551_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n568_), .A2(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT73), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n579_), .B(new_n552_), .C1(new_n576_), .C2(new_n551_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n581_), .A2(KEYINPUT37), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT37), .B1(new_n581_), .B2(new_n582_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT75), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n586_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT78), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n210_), .B(KEYINPUT74), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n298_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n594_), .B(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n264_), .B(new_n596_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n592_), .A3(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n598_), .A2(KEYINPUT79), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT79), .B1(new_n598_), .B2(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n583_), .A2(new_n584_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n548_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT99), .ZN(new_n607_));
  INV_X1    g406(.A(new_n536_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n607_), .A2(new_n291_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n609_), .A2(new_n610_), .A3(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n317_), .A2(new_n547_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n598_), .A2(new_n601_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n581_), .A2(new_n582_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT100), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n291_), .B1(new_n616_), .B2(new_n608_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n609_), .B2(KEYINPUT38), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n610_), .B1(new_n609_), .B2(KEYINPUT38), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n611_), .A2(new_n618_), .A3(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n543_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n292_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT39), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n607_), .A2(new_n292_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1325gat));
  INV_X1    g426(.A(G15gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n616_), .B2(new_n493_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n606_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n628_), .A3(new_n493_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n533_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n529_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n635_), .B1(new_n616_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT42), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  INV_X1    g441(.A(new_n604_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n612_), .A2(new_n643_), .A3(new_n614_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n608_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n547_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n614_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n581_), .A2(KEYINPUT37), .A3(new_n582_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(KEYINPUT43), .A3(new_n547_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n648_), .A2(new_n604_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(KEYINPUT44), .A3(new_n317_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(new_n608_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n648_), .A2(new_n604_), .A3(new_n317_), .A4(new_n653_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(G29gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n645_), .B1(new_n656_), .B2(new_n660_), .ZN(G1328gat));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n644_), .A2(new_n662_), .A3(new_n621_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT45), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n543_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n655_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT103), .B1(new_n666_), .B2(G36gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n668_), .B(new_n662_), .C1(new_n655_), .C2(new_n665_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT46), .B(new_n664_), .C1(new_n667_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  NAND2_X1  g473(.A1(new_n644_), .A2(new_n493_), .ZN(new_n675_));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n659_), .A2(G43gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n493_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n677_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1330gat));
  NAND3_X1  g485(.A1(new_n655_), .A2(new_n638_), .A3(new_n659_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G50gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT106), .ZN(new_n689_));
  INV_X1    g488(.A(new_n638_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(G50gat), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n644_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n689_), .A2(new_n693_), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n289_), .A2(new_n316_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n547_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n643_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n536_), .A4(new_n615_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n652_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n536_), .B1(new_n700_), .B2(KEYINPUT108), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(KEYINPUT108), .B2(new_n700_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n699_), .B1(new_n702_), .B2(new_n698_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n697_), .A2(new_n615_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n621_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT48), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n700_), .A2(new_n704_), .A3(new_n621_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1333gat));
  INV_X1    g508(.A(G71gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n705_), .B2(new_n493_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT49), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n700_), .A2(new_n710_), .A3(new_n493_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n705_), .A2(new_n638_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G78gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n717_), .A3(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n716_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n721_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n723_), .A2(KEYINPUT109), .A3(new_n719_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n715_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n690_), .A2(G78gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT111), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n700_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT109), .B1(new_n723_), .B2(new_n719_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n720_), .A2(new_n716_), .A3(new_n721_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(KEYINPUT50), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n725_), .A2(new_n728_), .A3(new_n731_), .ZN(G1335gat));
  AND4_X1   g531(.A1(new_n604_), .A2(new_n696_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n608_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n648_), .A2(new_n604_), .A3(new_n653_), .A4(new_n695_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n608_), .A2(G85gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT112), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n736_), .B2(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n733_), .B2(new_n621_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT113), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n621_), .A2(G92gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n736_), .B2(new_n742_), .ZN(G1337gat));
  INV_X1    g542(.A(new_n242_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n744_), .A3(new_n493_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G99gat), .B1(new_n735_), .B2(new_n492_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g547(.A1(new_n654_), .A2(KEYINPUT114), .A3(new_n638_), .A4(new_n695_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n735_), .B2(new_n690_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(G106gat), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT52), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n749_), .A2(new_n754_), .A3(new_n751_), .A4(G106gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n733_), .A2(new_n215_), .A3(new_n638_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  INV_X1    g562(.A(new_n316_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n605_), .A2(new_n763_), .A3(new_n764_), .A4(new_n289_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n650_), .A2(new_n643_), .A3(new_n651_), .A4(new_n289_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT54), .B1(new_n766_), .B2(new_n316_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n310_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n311_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n310_), .A2(new_n769_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n306_), .A2(new_n311_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n315_), .A3(new_n774_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n312_), .A2(new_n315_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT117), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n776_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n783_));
  NAND2_X1  g582(.A1(new_n271_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n267_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n249_), .A2(new_n272_), .A3(new_n262_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n785_), .A2(KEYINPUT55), .B1(new_n786_), .B2(new_n263_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n278_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n783_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n263_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n267_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT56), .B(new_n278_), .C1(new_n791_), .C2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n287_), .B(new_n782_), .C1(new_n789_), .C2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n278_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n280_), .B1(new_n802_), .B2(new_n795_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT58), .A3(new_n782_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n652_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n287_), .A2(new_n316_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n802_), .B2(new_n795_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n781_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n614_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n614_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT118), .A3(new_n813_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n799_), .A2(new_n652_), .A3(new_n817_), .A4(new_n804_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n806_), .A2(new_n815_), .A3(new_n816_), .A4(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n768_), .B1(new_n819_), .B2(new_n613_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n621_), .A2(new_n536_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n545_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n316_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT59), .B1(new_n820_), .B2(new_n822_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n805_), .A2(new_n814_), .A3(new_n810_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n604_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n765_), .A2(new_n767_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n545_), .A4(new_n821_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n825_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n316_), .A2(G113gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT120), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n824_), .B1(new_n832_), .B2(new_n834_), .ZN(G1340gat));
  INV_X1    g634(.A(new_n289_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n825_), .A2(new_n836_), .A3(new_n831_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT121), .B(G120gat), .Z(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n838_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n823_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(G1341gat));
  INV_X1    g642(.A(new_n613_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n825_), .A2(G127gat), .A3(new_n844_), .A4(new_n831_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n819_), .A2(new_n613_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n828_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n822_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n643_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n845_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n845_), .A2(new_n854_), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n832_), .A2(G134gat), .A3(new_n652_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n823_), .A2(new_n615_), .ZN(new_n858_));
  INV_X1    g657(.A(G134gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1343gat));
  INV_X1    g660(.A(new_n544_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n820_), .A2(new_n862_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(new_n821_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n316_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G141gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n327_), .A3(new_n316_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n836_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G148gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n328_), .A3(new_n836_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1345gat));
  NAND4_X1  g671(.A1(new_n847_), .A2(new_n643_), .A3(new_n544_), .A4(new_n821_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT123), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n863_), .A2(new_n875_), .A3(new_n643_), .A4(new_n821_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  NAND2_X1  g679(.A1(new_n864_), .A2(new_n615_), .ZN(new_n881_));
  INV_X1    g680(.A(G162gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n652_), .A2(G162gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT124), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n864_), .B2(new_n884_), .ZN(G1347gat));
  AND2_X1   g684(.A1(new_n829_), .A2(new_n545_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n608_), .A2(new_n543_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888_), .B2(new_n764_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n886_), .A2(new_n887_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n316_), .A3(new_n396_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT62), .B(G169gat), .C1(new_n888_), .C2(new_n764_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  NOR2_X1   g694(.A1(new_n820_), .A2(new_n638_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n608_), .A2(new_n543_), .A3(new_n492_), .ZN(new_n897_));
  AND4_X1   g696(.A1(G176gat), .A2(new_n896_), .A3(new_n836_), .A4(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n397_), .B1(new_n888_), .B2(new_n289_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT125), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n901_), .B(new_n397_), .C1(new_n888_), .C2(new_n289_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n898_), .B1(new_n900_), .B2(new_n902_), .ZN(G1349gat));
  INV_X1    g702(.A(new_n418_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n896_), .A2(new_n643_), .A3(new_n897_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n844_), .A2(new_n391_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n892_), .B2(new_n906_), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n892_), .A2(new_n392_), .A3(new_n615_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n652_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G190gat), .B1(new_n888_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n863_), .A2(new_n316_), .A3(new_n887_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n863_), .A2(new_n887_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT126), .B(G204gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n836_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n916_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n914_), .B2(new_n289_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1353gat));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  AND4_X1   g720(.A1(new_n844_), .A2(new_n847_), .A3(new_n544_), .A4(new_n887_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n921_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n925_));
  OAI211_X1 g724(.A(KEYINPUT127), .B(new_n923_), .C1(new_n914_), .C2(new_n613_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT63), .B(G211gat), .Z(new_n927_));
  AOI22_X1  g726(.A1(new_n925_), .A2(new_n926_), .B1(new_n922_), .B2(new_n927_), .ZN(G1354gat));
  INV_X1    g727(.A(G218gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n914_), .A2(new_n929_), .A3(new_n909_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n915_), .A2(new_n615_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(new_n931_), .ZN(G1355gat));
endmodule


