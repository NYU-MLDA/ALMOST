//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_;
  XNOR2_X1  g000(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT34), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT35), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G85gat), .B(G92gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT8), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n223_), .A2(KEYINPUT66), .A3(new_n219_), .A4(new_n218_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n216_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n210_), .B1(new_n225_), .B2(KEYINPUT67), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227_));
  AOI211_X1 g026(.A(new_n227_), .B(new_n216_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT68), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n222_), .A2(new_n224_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n227_), .B1(new_n230_), .B2(new_n216_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(KEYINPUT67), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .A4(new_n210_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n209_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(new_n213_), .B2(new_n215_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n211_), .A3(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(KEYINPUT70), .B(new_n235_), .C1(new_n230_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n222_), .A2(new_n224_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n244_), .A2(new_n211_), .A3(new_n236_), .A4(new_n240_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT70), .B1(new_n245_), .B2(new_n235_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n229_), .B(new_n234_), .C1(new_n243_), .C2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT10), .B(G99gat), .Z(new_n248_));
  INV_X1    g047(.A(G106gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n248_), .A2(new_n249_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n235_), .A2(new_n251_), .A3(KEYINPUT9), .ZN(new_n252_));
  INV_X1    g051(.A(G85gat), .ZN(new_n253_));
  INV_X1    g052(.A(G92gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT9), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n209_), .B2(KEYINPUT64), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n247_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G29gat), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G43gat), .B(G50gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT15), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n208_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n247_), .A2(new_n261_), .A3(new_n257_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n206_), .A2(new_n207_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n247_), .A2(KEYINPUT73), .A3(new_n261_), .A4(new_n257_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n263_), .A2(new_n266_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n264_), .A2(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n267_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n266_), .A2(KEYINPUT74), .A3(new_n267_), .A4(new_n268_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n258_), .A2(new_n262_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n258_), .A2(KEYINPUT72), .A3(new_n262_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(new_n275_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n270_), .B1(new_n280_), .B2(new_n208_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G190gat), .B(G218gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT75), .ZN(new_n283_));
  XOR2_X1   g082(.A(G134gat), .B(G162gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT36), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  AOI211_X1 g088(.A(new_n270_), .B(new_n289_), .C1(new_n280_), .C2(new_n208_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n203_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n208_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n289_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n269_), .A3(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(new_n202_), .C1(new_n281_), .C2(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT16), .ZN(new_n299_));
  XOR2_X1   g098(.A(G183gat), .B(G211gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT17), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT77), .Z(new_n304_));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305_));
  INV_X1    g104(.A(G1gat), .ZN(new_n306_));
  INV_X1    g105(.A(G8gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT14), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G8gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n315_));
  XOR2_X1   g114(.A(G71gat), .B(G78gat), .Z(new_n316_));
  OR2_X1    g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n316_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n313_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n304_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n320_), .B(KEYINPUT71), .Z(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(new_n313_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n313_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n302_), .A2(KEYINPUT17), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n303_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n297_), .A2(new_n328_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n247_), .A2(new_n257_), .A3(new_n323_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n320_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n247_), .B2(new_n257_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n323_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n258_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G230gat), .A2(G233gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n247_), .A2(new_n257_), .A3(new_n323_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G120gat), .B(G148gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT5), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G176gat), .B(G204gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n339_), .A2(new_n343_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT13), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(KEYINPUT13), .A3(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n311_), .B(new_n261_), .Z(new_n357_));
  NAND2_X1  g156(.A1(G229gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT78), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n262_), .A2(new_n311_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n311_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n261_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n364_), .A3(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G141gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G169gat), .B(G197gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n369_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n356_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT23), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  INV_X1    g177(.A(G176gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT24), .A3(new_n381_), .ZN(new_n382_));
  OR3_X1    g181(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n377_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n377_), .B1(G183gat), .B2(G190gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT81), .B(G176gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT22), .B(G169gat), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n390_), .A2(new_n391_), .B1(G169gat), .B2(G176gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G197gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(G204gat), .ZN(new_n396_));
  INV_X1    g195(.A(G204gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(G197gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT21), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n395_), .B2(G204gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n402_), .B(new_n403_), .C1(G197gat), .C2(new_n397_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n399_), .B(new_n400_), .C1(new_n404_), .C2(KEYINPUT21), .ZN(new_n405_));
  INV_X1    g204(.A(new_n400_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(KEYINPUT21), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n394_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT19), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT94), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT26), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT79), .B1(new_n414_), .B2(G190gat), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n415_), .B(new_n386_), .C1(new_n385_), .C2(KEYINPUT79), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT80), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n414_), .A2(G190gat), .ZN(new_n419_));
  INV_X1    g218(.A(G190gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(KEYINPUT26), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n415_), .A4(new_n386_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n384_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n393_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT82), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n428_), .A3(new_n393_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n413_), .B1(new_n430_), .B2(new_n408_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n425_), .A2(new_n428_), .A3(new_n393_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n428_), .B1(new_n425_), .B2(new_n393_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n413_), .B(new_n408_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n412_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n411_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n405_), .A2(new_n407_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n384_), .A2(new_n387_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n394_), .A2(KEYINPUT93), .A3(new_n408_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n438_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n427_), .A2(new_n429_), .A3(new_n440_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n437_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n436_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT96), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n452_), .B(new_n453_), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n432_), .A2(new_n433_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT94), .B1(new_n456_), .B2(new_n440_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n434_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n446_), .B1(new_n458_), .B2(new_n412_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT27), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n444_), .A2(new_n437_), .A3(new_n445_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n409_), .A2(KEYINPUT98), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT98), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(KEYINPUT20), .C1(new_n394_), .C2(new_n408_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n457_), .B2(new_n434_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n464_), .B1(new_n469_), .B2(new_n437_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n454_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n463_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n462_), .A2(new_n463_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT0), .B(G57gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n478_));
  INV_X1    g277(.A(G141gat), .ZN(new_n479_));
  INV_X1    g278(.A(G148gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT3), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487_));
  OR2_X1    g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G141gat), .B(G148gat), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(KEYINPUT1), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n488_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n487_), .A2(KEYINPUT1), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G127gat), .B(G134gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G113gat), .B(G120gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G120gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n489_), .A2(new_n494_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(KEYINPUT84), .A3(new_n501_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G225gat), .A2(G233gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n499_), .A2(KEYINPUT84), .A3(new_n501_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT84), .B1(new_n499_), .B2(new_n501_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT4), .B1(new_n516_), .B2(new_n506_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n477_), .B(new_n511_), .C1(new_n518_), .C2(new_n510_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n477_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n513_), .A2(new_n517_), .A3(new_n510_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n511_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n473_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n456_), .A2(KEYINPUT30), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n430_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n527_), .A2(new_n529_), .A3(KEYINPUT83), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT83), .B1(new_n527_), .B2(new_n529_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G43gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G227gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(G15gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n534_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n530_), .A2(new_n531_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n539_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n516_), .B(KEYINPUT31), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT85), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n542_), .A2(KEYINPUT85), .ZN(new_n545_));
  OR3_X1    g344(.A1(new_n540_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n440_), .B2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT90), .B(new_n408_), .C1(new_n495_), .C2(new_n548_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT87), .B(G228gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT88), .B(G233gat), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n550_), .B(new_n551_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n440_), .A2(new_n549_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n553_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(KEYINPUT90), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G78gat), .B(G106gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n495_), .A2(new_n548_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT28), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G22gat), .B(G50gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n560_), .B1(new_n558_), .B2(KEYINPUT91), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n554_), .A2(new_n567_), .A3(new_n557_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n566_), .A2(KEYINPUT92), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT92), .B1(new_n566_), .B2(new_n568_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n561_), .B(new_n565_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n545_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n558_), .B(new_n560_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n565_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n565_), .A2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n573_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n546_), .A2(new_n571_), .A3(new_n572_), .A4(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n526_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n460_), .A2(KEYINPUT32), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n465_), .A2(new_n467_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n411_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n581_), .B1(new_n584_), .B2(new_n464_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n436_), .A2(new_n581_), .A3(new_n447_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n524_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n580_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n459_), .A2(new_n581_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n581_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n470_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n591_), .A3(KEYINPUT99), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n477_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n518_), .B2(new_n510_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n523_), .A2(KEYINPUT97), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(KEYINPUT33), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n523_), .A2(KEYINPUT97), .A3(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n596_), .A2(new_n455_), .A3(new_n461_), .A4(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n571_), .A2(new_n577_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n524_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n473_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n546_), .A2(new_n572_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n579_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n375_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n329_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT100), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n306_), .A3(new_n524_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT101), .B1(new_n288_), .B2(new_n290_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n294_), .B(new_n617_), .C1(new_n281_), .C2(new_n287_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n600_), .A2(new_n601_), .B1(new_n603_), .B2(new_n473_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n606_), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n620_), .A2(new_n621_), .B1(new_n578_), .B2(new_n526_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT102), .ZN(new_n624_));
  INV_X1    g423(.A(new_n328_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n374_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n624_), .A2(KEYINPUT103), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT103), .B1(new_n624_), .B2(new_n627_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n524_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n631_), .A2(KEYINPUT104), .A3(G1gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT104), .B1(new_n631_), .B2(G1gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n615_), .B1(new_n632_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n473_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n610_), .A2(new_n307_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n624_), .A2(new_n635_), .A3(new_n627_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n624_), .A2(new_n639_), .A3(new_n635_), .A4(new_n627_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G8gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n637_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n638_), .A2(new_n639_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(new_n642_), .A3(KEYINPUT39), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n636_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT40), .B(new_n636_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  NAND3_X1  g450(.A1(new_n610_), .A2(new_n536_), .A3(new_n621_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n621_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n653_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n653_), .B2(G15gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n652_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT107), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n658_), .B(new_n652_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n601_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n610_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n630_), .A2(new_n662_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G22gat), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT42), .B(new_n661_), .C1(new_n630_), .C2(new_n662_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(G1327gat));
  OAI21_X1  g467(.A(KEYINPUT43), .B1(new_n607_), .B2(new_n296_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n622_), .A2(new_n670_), .A3(new_n295_), .A4(new_n291_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n374_), .A2(new_n328_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n676_), .B(new_n673_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n525_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n619_), .A2(new_n625_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n608_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n608_), .A3(KEYINPUT108), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n686_), .A2(G29gat), .A3(new_n525_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n680_), .A2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n672_), .A2(new_n674_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n676_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n674_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n635_), .A4(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n678_), .B2(new_n635_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n473_), .A2(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n684_), .A2(new_n685_), .A3(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n691_), .A2(new_n635_), .A3(new_n693_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT109), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(KEYINPUT110), .A3(G36gat), .A4(new_n694_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n697_), .A2(new_n702_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n706_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(G36gat), .A3(new_n694_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n701_), .B1(new_n712_), .B2(new_n689_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n713_), .A2(new_n707_), .A3(new_n708_), .A4(new_n705_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1329gat));
  OAI21_X1  g514(.A(G43gat), .B1(new_n679_), .B2(new_n606_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n621_), .A2(new_n533_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n686_), .B2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n679_), .B2(new_n601_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n601_), .A2(G50gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT113), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n686_), .B2(new_n722_), .ZN(G1331gat));
  INV_X1    g522(.A(new_n356_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n372_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n624_), .A2(new_n625_), .A3(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(G57gat), .A3(new_n524_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n607_), .A2(new_n372_), .A3(new_n724_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n329_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n525_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n727_), .A2(new_n728_), .B1(G57gat), .B2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n728_), .B2(new_n727_), .ZN(G1332gat));
  INV_X1    g532(.A(G64gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n726_), .B2(new_n635_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT48), .Z(new_n736_));
  INV_X1    g535(.A(new_n730_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n734_), .A3(new_n635_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n726_), .B2(new_n621_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n621_), .A2(new_n740_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT116), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n730_), .B2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n726_), .B2(new_n662_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n737_), .A2(new_n747_), .A3(new_n662_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1335gat));
  AND2_X1   g551(.A1(new_n729_), .A2(new_n681_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n253_), .A3(new_n524_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n672_), .A2(new_n328_), .A3(new_n725_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n524_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(new_n253_), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n254_), .A3(new_n635_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n755_), .A2(new_n635_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n254_), .ZN(G1337gat));
  INV_X1    g559(.A(G99gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n755_), .B2(new_n621_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT118), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n621_), .A2(new_n248_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n753_), .A2(new_n764_), .B1(KEYINPUT119), .B2(KEYINPUT51), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n766_), .B(new_n767_), .Z(G1338gat));
  AOI21_X1  g567(.A(new_n249_), .B1(new_n755_), .B2(new_n662_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT52), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n753_), .A2(new_n249_), .A3(new_n662_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g572(.A(new_n578_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n635_), .A2(new_n525_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n357_), .A2(new_n358_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n362_), .A2(new_n364_), .A3(new_n359_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n369_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n370_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n352_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n338_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n339_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n332_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n258_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n340_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT12), .B1(new_n258_), .B2(new_n335_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n782_), .A4(new_n342_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n348_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n792_), .B(new_n350_), .C1(new_n783_), .C2(new_n789_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n791_), .A2(new_n793_), .A3(KEYINPUT121), .ZN(new_n794_));
  NOR4_X1   g593(.A1(new_n787_), .A2(new_n330_), .A3(new_n342_), .A4(new_n333_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n342_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(KEYINPUT55), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n348_), .B1(new_n797_), .B2(new_n788_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT121), .A3(new_n792_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n372_), .A2(new_n351_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n780_), .B1(new_n794_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n619_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n792_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n348_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n779_), .A2(new_n351_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT58), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n812_), .B(new_n809_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n804_), .A2(new_n805_), .B1(new_n814_), .B2(new_n297_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n803_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n625_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n373_), .A2(new_n625_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT120), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n296_), .A2(new_n724_), .A3(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n774_), .B(new_n775_), .C1(new_n817_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n372_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n806_), .A2(new_n829_), .A3(new_n807_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n800_), .B1(new_n791_), .B2(KEYINPUT121), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n830_), .A2(new_n831_), .B1(new_n352_), .B2(new_n779_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n616_), .A2(new_n618_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n805_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n808_), .A2(new_n810_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n812_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n810_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n297_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n816_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n328_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n821_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .A3(new_n774_), .A4(new_n775_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n373_), .B1(new_n828_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n826_), .B1(new_n843_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n845_));
  AOI21_X1  g644(.A(G120gat), .B1(new_n356_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT122), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n845_), .B2(G120gat), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n824_), .B(new_n847_), .C1(new_n846_), .C2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n724_), .B1(new_n828_), .B2(new_n842_), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n824_), .A2(new_n854_), .A3(new_n625_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n328_), .B1(new_n828_), .B2(new_n842_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n854_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT123), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n855_), .C1(new_n856_), .C2(new_n854_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n824_), .A2(new_n862_), .A3(new_n833_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n296_), .B1(new_n828_), .B2(new_n842_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1343gat));
  AND2_X1   g664(.A1(new_n841_), .A2(new_n775_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n621_), .A2(new_n601_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n373_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n479_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n724_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n480_), .ZN(G1345gat));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n868_), .B2(new_n328_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n866_), .A2(KEYINPUT124), .A3(new_n625_), .A4(new_n867_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n868_), .B2(new_n296_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n619_), .A2(G162gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n868_), .B2(new_n881_), .ZN(G1347gat));
  AOI211_X1 g681(.A(new_n524_), .B(new_n473_), .C1(new_n840_), .C2(new_n821_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n774_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n373_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n885_), .A2(new_n378_), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n885_), .B2(new_n378_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n391_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1348gat));
  NAND3_X1  g689(.A1(new_n883_), .A2(new_n774_), .A3(new_n356_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n379_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n390_), .B2(new_n891_), .ZN(G1349gat));
  NOR2_X1   g692(.A1(new_n884_), .A2(new_n328_), .ZN(new_n894_));
  MUX2_X1   g693(.A(G183gat), .B(new_n386_), .S(new_n894_), .Z(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n884_), .B2(new_n296_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n833_), .A2(new_n385_), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT126), .Z(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n884_), .B2(new_n898_), .ZN(G1351gat));
  NAND2_X1  g698(.A1(new_n883_), .A2(new_n867_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n373_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n395_), .ZN(G1352gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n724_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n397_), .ZN(G1353gat));
  OAI22_X1  g703(.A1(new_n900_), .A2(new_n328_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n883_), .A2(new_n625_), .A3(new_n867_), .A4(new_n907_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n905_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n906_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1354gat));
  OAI21_X1  g710(.A(G218gat), .B1(new_n900_), .B2(new_n296_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n619_), .A2(G218gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n900_), .B2(new_n913_), .ZN(G1355gat));
endmodule


