//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT89), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT88), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n208_), .B2(KEYINPUT1), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT90), .B(KEYINPUT2), .Z(new_n218_));
  NOR2_X1   g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT91), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  OAI22_X1  g021(.A1(new_n215_), .A2(new_n221_), .B1(new_n212_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n221_), .B2(new_n215_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n208_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n204_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n217_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT84), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT85), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n232_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n228_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n235_), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n217_), .B1(new_n238_), .B2(new_n233_), .C1(new_n225_), .C2(new_n227_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n203_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT4), .B1(new_n228_), .B2(new_n236_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n240_), .B1(new_n244_), .B2(new_n203_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n245_), .B(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT31), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(KEYINPUT31), .A3(new_n253_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT83), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G15gat), .B(G43gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT82), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT30), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G169gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT80), .B(G183gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(G190gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n264_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(KEYINPUT25), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT81), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(G169gat), .B2(G176gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n279_), .B(new_n266_), .C1(KEYINPUT24), .C2(new_n276_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n270_), .B1(new_n274_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(G71gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G99gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n281_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n261_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT83), .A4(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n262_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n286_), .B1(new_n262_), .B2(new_n288_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n251_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT96), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n294_), .A2(new_n273_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(new_n280_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n264_), .B1(new_n267_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300_));
  AND2_X1   g099(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(KEYINPUT20), .C1(new_n307_), .C2(new_n281_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT101), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n307_), .B1(new_n299_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n313_), .B2(new_n299_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n281_), .A2(new_n307_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT97), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(KEYINPUT97), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n315_), .A2(KEYINPUT20), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n312_), .B1(new_n319_), .B2(new_n311_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G8gat), .B(G36gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G64gat), .B(G92gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n320_), .A2(KEYINPUT102), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n309_), .A2(new_n311_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n296_), .A2(new_n298_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n311_), .B1(new_n328_), .B2(new_n306_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n329_), .A2(new_n318_), .A3(KEYINPUT20), .A4(new_n317_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n325_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT27), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n326_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT102), .B1(new_n320_), .B2(new_n325_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n325_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n334_), .A2(new_n335_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G50gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(new_n217_), .C1(new_n225_), .C2(new_n227_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G22gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n345_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n342_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G22gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(G50gat), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n306_), .B1(new_n228_), .B2(KEYINPUT29), .ZN(new_n357_));
  OAI21_X1  g156(.A(G233gat), .B1(KEYINPUT92), .B2(G228gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(KEYINPUT92), .B2(G228gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n306_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n357_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT94), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT95), .B1(new_n356_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n363_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n362_), .A2(new_n363_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT94), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n355_), .A4(new_n351_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n365_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n369_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n291_), .B(new_n341_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n320_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(KEYINPUT100), .Z(new_n380_));
  NAND2_X1  g179(.A1(new_n331_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n244_), .A2(new_n203_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n240_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n249_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n245_), .A2(new_n250_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n379_), .B(new_n381_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n237_), .A2(new_n239_), .A3(new_n203_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n250_), .B(new_n388_), .C1(new_n244_), .C2(new_n203_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n332_), .A3(new_n338_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(new_n391_), .A3(new_n249_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT33), .B1(new_n245_), .B2(new_n250_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n387_), .B1(new_n394_), .B2(KEYINPUT99), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT99), .ZN(new_n396_));
  AOI211_X1 g195(.A(new_n396_), .B(new_n390_), .C1(new_n393_), .C2(new_n392_), .ZN(new_n397_));
  OAI22_X1  g196(.A1(new_n395_), .A2(new_n397_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n365_), .A2(new_n373_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n369_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n251_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n365_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n401_), .A2(new_n341_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n289_), .A2(new_n290_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n377_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G64gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G57gat), .ZN(new_n411_));
  INV_X1    g210(.A(G57gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G64gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT11), .ZN(new_n414_));
  INV_X1    g213(.A(G78gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G71gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n283_), .A2(G78gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n414_), .A2(new_n418_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G57gat), .B(G64gat), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n421_), .A2(KEYINPUT11), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT12), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n429_));
  INV_X1    g228(.A(G99gat), .ZN(new_n430_));
  INV_X1    g229(.A(G106gat), .ZN(new_n431_));
  OAI22_X1  g230(.A1(new_n427_), .A2(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n438_));
  AND2_X1   g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n432_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT8), .ZN(new_n442_));
  OR2_X1    g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n441_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G92gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT9), .ZN(new_n451_));
  AND2_X1   g250(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n431_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n443_), .A2(KEYINPUT9), .A3(new_n444_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n439_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(KEYINPUT66), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n432_), .A2(new_n440_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n449_), .A2(KEYINPUT67), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n463_), .A2(new_n467_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n433_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n460_), .A2(new_n461_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT8), .B1(new_n475_), .B2(new_n445_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n441_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n470_), .B1(new_n471_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n425_), .B1(new_n469_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G230gat), .A2(G233gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n465_), .A2(new_n466_), .ZN(new_n482_));
  AOI211_X1 g281(.A(new_n482_), .B(new_n423_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n423_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n483_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n481_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT68), .ZN(new_n490_));
  INV_X1    g289(.A(new_n423_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n478_), .B2(new_n484_), .ZN(new_n492_));
  OAI211_X1 g291(.A(G230gat), .B(G233gat), .C1(new_n492_), .C2(new_n483_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n480_), .A2(new_n494_), .A3(new_n488_), .A4(new_n481_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G120gat), .B(G148gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(G176gat), .B(G204gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n490_), .A2(new_n493_), .A3(new_n495_), .A4(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n502_), .A2(KEYINPUT13), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT13), .B1(new_n502_), .B2(new_n504_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G1gat), .ZN(new_n509_));
  INV_X1    g308(.A(G8gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT74), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT74), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G1gat), .B(G8gat), .Z(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  XNOR2_X1  g316(.A(G29gat), .B(G36gat), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT70), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT70), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n524_), .A2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT15), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n532_), .B2(new_n517_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT78), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n517_), .B(new_n526_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n534_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n533_), .A2(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT79), .ZN(new_n540_));
  XOR2_X1   g339(.A(G169gat), .B(G197gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n538_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n508_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n409_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT104), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT72), .ZN(new_n549_));
  XOR2_X1   g348(.A(G134gat), .B(G162gat), .Z(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  OAI21_X1  g350(.A(new_n532_), .B1(new_n469_), .B2(new_n479_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n485_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n528_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n552_), .A2(KEYINPUT71), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT67), .B1(new_n449_), .B2(new_n468_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n471_), .A2(new_n478_), .A3(new_n470_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n564_), .A2(new_n565_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n568_), .A3(new_n554_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n562_), .B1(new_n569_), .B2(new_n558_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n551_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n551_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n566_), .A2(new_n567_), .B1(new_n528_), .B2(new_n553_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n557_), .B1(new_n576_), .B2(new_n563_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT73), .B1(new_n577_), .B2(new_n562_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n554_), .B1(new_n552_), .B2(KEYINPUT71), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n566_), .A2(new_n567_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n558_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n571_), .B1(new_n583_), .B2(new_n561_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n578_), .B(new_n574_), .C1(new_n584_), .C2(new_n573_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(KEYINPUT37), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  INV_X1    g386(.A(new_n585_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n578_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n423_), .B(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT75), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n517_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT77), .ZN(new_n597_));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT17), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n597_), .B(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n596_), .A2(KEYINPUT17), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n592_), .A2(new_n606_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n546_), .A2(new_n547_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n547_), .B1(new_n546_), .B2(new_n607_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n509_), .A3(new_n251_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n610_), .A2(KEYINPUT38), .A3(new_n509_), .A4(new_n251_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n580_), .A2(new_n585_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n606_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n409_), .A2(new_n545_), .A3(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n402_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n613_), .A2(new_n614_), .A3(new_n620_), .ZN(G1324gat));
  INV_X1    g420(.A(new_n341_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n608_), .A2(new_n510_), .A3(new_n622_), .A4(new_n609_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G8gat), .B1(new_n619_), .B2(new_n341_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(G8gat), .C1(new_n619_), .C2(new_n341_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n610_), .A2(new_n632_), .A3(new_n406_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G15gat), .B1(new_n619_), .B2(new_n407_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  NAND2_X1  g436(.A1(new_n401_), .A2(new_n403_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n610_), .A2(new_n347_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G22gat), .B1(new_n619_), .B2(new_n638_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT42), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT43), .B1(new_n408_), .B2(new_n592_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n406_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n646_), .B(new_n591_), .C1(new_n647_), .C2(new_n377_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n545_), .A2(new_n617_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n251_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G29gat), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n615_), .A2(new_n606_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n409_), .A2(new_n658_), .A3(new_n545_), .A4(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n545_), .B(new_n659_), .C1(new_n647_), .C2(new_n377_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT105), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n663_), .A2(G29gat), .A3(new_n402_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n644_), .B1(new_n657_), .B2(new_n665_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT106), .B(new_n664_), .C1(new_n656_), .C2(G29gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n660_), .A2(new_n669_), .A3(new_n622_), .A4(new_n662_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT45), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n649_), .B2(new_n651_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n653_), .B(new_n650_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n341_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n669_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n671_), .B(KEYINPUT46), .C1(new_n669_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  AND2_X1   g478(.A1(new_n660_), .A2(new_n662_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G43gat), .B1(new_n680_), .B2(new_n406_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n672_), .A2(new_n673_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n406_), .A2(G43gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1330gat));
  NAND3_X1  g485(.A1(new_n680_), .A2(new_n342_), .A3(new_n639_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n682_), .A2(new_n688_), .A3(new_n639_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n682_), .B2(new_n639_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NOR3_X1   g491(.A1(new_n408_), .A2(new_n543_), .A3(new_n507_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n618_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n402_), .ZN(new_n695_));
  NOR4_X1   g494(.A1(new_n408_), .A2(new_n543_), .A3(new_n507_), .A4(new_n607_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n412_), .A3(new_n251_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1332gat));
  NAND3_X1  g497(.A1(new_n696_), .A2(new_n410_), .A3(new_n622_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n694_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n622_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(G64gat), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n701_), .B2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n699_), .B1(new_n704_), .B2(new_n705_), .ZN(G1333gat));
  NAND3_X1  g505(.A1(new_n696_), .A2(new_n283_), .A3(new_n406_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n700_), .A2(new_n406_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(G71gat), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n708_), .B2(G71gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1334gat));
  NAND3_X1  g512(.A1(new_n696_), .A2(new_n415_), .A3(new_n639_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n700_), .A2(new_n639_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(G78gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n715_), .B2(G78gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(G1335gat));
  NAND2_X1  g519(.A1(new_n693_), .A2(new_n659_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n251_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n617_), .A2(new_n508_), .A3(new_n544_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT109), .Z(new_n726_));
  NOR2_X1   g525(.A1(new_n452_), .A2(new_n453_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n402_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n726_), .B2(new_n728_), .ZN(G1336gat));
  OAI21_X1  g528(.A(new_n450_), .B1(new_n721_), .B2(new_n341_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT110), .Z(new_n731_));
  NOR2_X1   g530(.A1(new_n341_), .A2(new_n450_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n726_), .B2(new_n732_), .ZN(G1337gat));
  AND2_X1   g532(.A1(new_n725_), .A2(new_n406_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n406_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n734_), .A2(new_n430_), .B1(new_n721_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n736_), .B(new_n737_), .Z(G1338gat));
  NAND3_X1  g537(.A1(new_n722_), .A2(new_n431_), .A3(new_n639_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n725_), .A2(new_n639_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G106gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT52), .B(new_n431_), .C1(new_n725_), .C2(new_n639_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n739_), .B(new_n745_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1339gat));
  NAND4_X1  g548(.A1(new_n638_), .A2(new_n251_), .A3(new_n341_), .A4(new_n406_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n542_), .B1(new_n536_), .B2(new_n535_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n535_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n533_), .A2(new_n753_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n538_), .A2(new_n542_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n504_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n490_), .A2(new_n757_), .A3(new_n495_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n424_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n478_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n492_), .B2(KEYINPUT12), .ZN(new_n761_));
  OAI211_X1 g560(.A(G230gat), .B(G233gat), .C1(new_n759_), .C2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n480_), .A2(KEYINPUT55), .A3(new_n488_), .A4(new_n481_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n758_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n501_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n767_), .B(new_n503_), .C1(new_n758_), .C2(new_n764_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n756_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT113), .B(new_n756_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n591_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT114), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n591_), .A3(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n769_), .A2(new_n772_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n766_), .A2(new_n768_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n543_), .A2(new_n504_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n502_), .A2(new_n504_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(new_n755_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n615_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT57), .B(new_n615_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n606_), .B1(new_n780_), .B2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n508_), .A2(new_n543_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n592_), .A2(new_n606_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n751_), .B1(new_n792_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT115), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n794_), .B(KEYINPUT54), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n778_), .A2(new_n779_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n790_), .B1(new_n800_), .B2(new_n776_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n801_), .B2(new_n606_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n751_), .ZN(new_n804_));
  INV_X1    g603(.A(G113gat), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n798_), .A2(new_n804_), .A3(new_n805_), .A4(new_n543_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n792_), .B2(new_n796_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n797_), .A3(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n802_), .B(new_n751_), .C1(KEYINPUT116), .C2(KEYINPUT59), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n544_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n811_), .B2(new_n805_), .ZN(G1340gat));
  NOR2_X1   g611(.A1(new_n507_), .A2(G120gat), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n798_), .B(new_n804_), .C1(KEYINPUT60), .C2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n507_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT117), .B(new_n507_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G120gat), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n814_), .A2(KEYINPUT60), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1341gat));
  INV_X1    g620(.A(G127gat), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n798_), .A2(new_n804_), .A3(new_n822_), .A4(new_n606_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n617_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n822_), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n798_), .A2(new_n804_), .A3(new_n826_), .A4(new_n616_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n592_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n826_), .ZN(G1343gat));
  NOR2_X1   g628(.A1(new_n792_), .A2(new_n796_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n407_), .A2(new_n341_), .A3(new_n251_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n830_), .A2(new_n638_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n543_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT118), .B(G141gat), .Z(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(G1344gat));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n508_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g636(.A1(new_n832_), .A2(new_n606_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT61), .B(G155gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1346gat));
  AOI21_X1  g639(.A(G162gat), .B1(new_n832_), .B2(new_n616_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n591_), .A2(G162gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT119), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n832_), .B2(new_n843_), .ZN(G1347gat));
  XNOR2_X1  g643(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n830_), .A2(new_n341_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n638_), .A2(new_n291_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n543_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n848_), .B2(KEYINPUT22), .ZN(new_n849_));
  OAI21_X1  g648(.A(G169gat), .B1(new_n848_), .B2(new_n845_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G169gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n849_), .ZN(G1348gat));
  NAND2_X1  g652(.A1(new_n846_), .A2(new_n847_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n508_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g656(.A(new_n268_), .B1(new_n854_), .B2(new_n617_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n846_), .A2(new_n294_), .A3(new_n606_), .A4(new_n847_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1350gat));
  NAND3_X1  g662(.A1(new_n855_), .A2(new_n273_), .A3(new_n616_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G190gat), .B1(new_n854_), .B2(new_n592_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(G1351gat));
  NOR3_X1   g667(.A1(new_n638_), .A2(new_n251_), .A3(new_n406_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n846_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n543_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g672(.A1(new_n870_), .A2(new_n507_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT123), .B(G204gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1353gat));
  NAND2_X1  g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n878_));
  INV_X1    g677(.A(G211gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(KEYINPUT124), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n871_), .A2(new_n606_), .A3(new_n877_), .A4(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n879_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1354gat));
  XNOR2_X1  g682(.A(KEYINPUT126), .B(G218gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n592_), .A2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT127), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n870_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n846_), .A2(new_n616_), .A3(new_n869_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT125), .Z(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n889_), .B2(new_n884_), .ZN(G1355gat));
endmodule


