//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT66), .B(G85gat), .Z(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n204_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT10), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT10), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(KEYINPUT10), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT64), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  AOI211_X1 g023(.A(new_n224_), .B(G106gat), .C1(new_n217_), .C2(new_n220_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n211_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT67), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n215_), .A2(new_n222_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT7), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n209_), .B(KEYINPUT6), .Z(new_n230_));
  OAI21_X1  g029(.A(new_n203_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n211_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G78gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n241_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n227_), .A2(new_n232_), .A3(new_n243_), .A4(new_n234_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(KEYINPUT12), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT12), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n235_), .A2(new_n246_), .A3(new_n241_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(KEYINPUT68), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n255_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n256_), .B2(new_n251_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G120gat), .B(G148gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT5), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G176gat), .ZN(new_n261_));
  INV_X1    g060(.A(G204gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n202_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  AOI211_X1 g064(.A(KEYINPUT69), .B(new_n265_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT13), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n256_), .A2(new_n251_), .A3(new_n263_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT68), .B1(new_n250_), .B2(new_n252_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n256_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n263_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT69), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n258_), .A2(new_n202_), .A3(new_n263_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n270_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT13), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G22gat), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  INV_X1    g080(.A(G8gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G1gat), .B(G8gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n241_), .B(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(G231gat), .A2(G233gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G155gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT16), .ZN(new_n291_));
  INV_X1    g090(.A(G183gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(G211gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT17), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n287_), .A2(new_n288_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT76), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n294_), .A2(new_n295_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  INV_X1    g100(.A(KEYINPUT15), .ZN(new_n302_));
  INV_X1    g101(.A(G29gat), .ZN(new_n303_));
  INV_X1    g102(.A(G36gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G29gat), .A2(G36gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n306_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n310_));
  OAI21_X1  g109(.A(G43gat), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n310_), .ZN(new_n312_));
  INV_X1    g111(.A(G43gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n308_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n314_), .A3(G50gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(G50gat), .B1(new_n311_), .B2(new_n314_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n302_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n311_), .A2(new_n314_), .ZN(new_n319_));
  INV_X1    g118(.A(G50gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(KEYINPUT15), .A3(new_n315_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n235_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT71), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G232gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT34), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(KEYINPUT35), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n315_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n235_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n324_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT35), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n324_), .B2(KEYINPUT71), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(new_n327_), .A3(new_n324_), .A4(new_n330_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n327_), .A2(KEYINPUT35), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G190gat), .B(G218gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT72), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G134gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G162gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n341_), .B(KEYINPUT36), .Z(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT37), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n337_), .A2(KEYINPUT74), .ZN(new_n347_));
  INV_X1    g146(.A(new_n344_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n332_), .A2(new_n335_), .A3(new_n349_), .A4(new_n336_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n343_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n301_), .B1(new_n346_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n279_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT77), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT77), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n366_));
  AND2_X1   g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT23), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n365_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT83), .B1(new_n366_), .B2(new_n367_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT84), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376_));
  OAI221_X1 g175(.A(new_n376_), .B1(G183gat), .B2(G190gat), .C1(new_n371_), .C2(new_n372_), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT22), .B1(new_n378_), .B2(KEYINPUT80), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(KEYINPUT81), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(KEYINPUT81), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n385_), .A2(KEYINPUT82), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n375_), .A2(new_n377_), .A3(new_n388_), .A4(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT78), .Z(new_n394_));
  OR2_X1    g193(.A1(new_n394_), .A2(KEYINPUT24), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n367_), .A2(new_n369_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n395_), .A2(new_n397_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n392_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n262_), .B2(G197gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(KEYINPUT21), .A3(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G197gat), .B(G204gat), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n406_), .A2(KEYINPUT21), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n406_), .A2(KEYINPUT21), .A3(new_n410_), .A4(new_n408_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n364_), .B1(new_n403_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n397_), .B1(G183gat), .B2(G190gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT22), .B(G169gat), .Z(new_n418_));
  OAI211_X1 g217(.A(new_n417_), .B(new_n386_), .C1(G176gat), .C2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n394_), .A2(new_n386_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n393_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n421_), .B(new_n400_), .C1(new_n422_), .C2(new_n420_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(new_n373_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n415_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n416_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT19), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n392_), .A2(new_n432_), .A3(new_n402_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n415_), .A2(new_n424_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n433_), .A2(KEYINPUT20), .A3(new_n434_), .A4(new_n429_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n363_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n429_), .B1(new_n416_), .B2(new_n426_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n363_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n358_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G141gat), .A2(G148gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT2), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n444_), .A2(KEYINPUT88), .A3(new_n445_), .A4(new_n447_), .ZN(new_n452_));
  OR2_X1    g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n451_), .A2(KEYINPUT1), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(KEYINPUT1), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G127gat), .B(G134gat), .ZN(new_n460_));
  INV_X1    g259(.A(G113gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G120gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n458_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n452_), .A2(new_n453_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n448_), .A2(new_n449_), .B1(G155gat), .B2(G162gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n463_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n464_), .A2(new_n470_), .A3(KEYINPUT4), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR3_X1    g272(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT4), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n464_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G85gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n475_), .A2(new_n482_), .A3(new_n476_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n432_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n488_), .A2(new_n425_), .A3(new_n364_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n435_), .B1(new_n489_), .B2(new_n429_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n439_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n433_), .A2(KEYINPUT20), .A3(new_n434_), .A4(new_n430_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n489_), .B2(new_n430_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n363_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n494_), .A3(KEYINPUT27), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n441_), .A2(new_n487_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G22gat), .B(G50gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT28), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n498_), .B1(new_n468_), .B2(new_n499_), .ZN(new_n500_));
  AND4_X1   g299(.A1(new_n498_), .A2(new_n454_), .A3(new_n499_), .A4(new_n458_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT89), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G228gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT28), .B1(new_n459_), .B2(KEYINPUT29), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n468_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n502_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n504_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n497_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT90), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n415_), .B(new_n512_), .C1(new_n499_), .C2(new_n468_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G78gat), .B(G106gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NOR3_X1   g314(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT89), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n506_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n503_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n502_), .A2(new_n508_), .A3(new_n504_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n497_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n511_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n515_), .B1(new_n511_), .B2(new_n521_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n392_), .A2(new_n526_), .A3(new_n402_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n525_), .B(new_n463_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n469_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n403_), .A2(KEYINPUT30), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(KEYINPUT85), .A3(new_n527_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n535_));
  XOR2_X1   g334(.A(G71gat), .B(G99gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G43gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G227gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n534_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n535_), .B1(new_n534_), .B2(new_n540_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n530_), .B(new_n532_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n532_), .A2(new_n530_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n540_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT31), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n543_), .A2(new_n548_), .A3(KEYINPUT86), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n496_), .A2(new_n524_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n439_), .A2(KEYINPUT32), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n493_), .A2(KEYINPUT98), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT98), .B1(new_n493_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n486_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n554_), .B(KEYINPUT96), .Z(new_n558_));
  AND3_X1   g357(.A1(new_n490_), .A2(KEYINPUT97), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT97), .B1(new_n490_), .B2(new_n558_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT99), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n493_), .A2(new_n554_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n493_), .A2(KEYINPUT98), .A3(new_n554_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n490_), .A2(new_n558_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n490_), .A2(KEYINPUT97), .A3(new_n558_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n567_), .A2(new_n572_), .A3(new_n573_), .A4(new_n486_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n515_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n509_), .A2(new_n510_), .A3(new_n497_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n520_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n575_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n511_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n436_), .A2(new_n440_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n464_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n581_), .A2(new_n483_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n485_), .A2(KEYINPUT33), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n475_), .A2(new_n585_), .A3(new_n482_), .A4(new_n476_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n583_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n578_), .A2(new_n579_), .B1(new_n580_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n562_), .A2(new_n574_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n553_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n524_), .A2(new_n549_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n496_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n323_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(new_n286_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n321_), .A2(new_n286_), .A3(new_n315_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n329_), .B(new_n286_), .Z(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n378_), .ZN(new_n604_));
  INV_X1    g403(.A(G197gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n594_), .A2(KEYINPUT100), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n553_), .A2(new_n589_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(new_n611_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n356_), .A2(new_n357_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n281_), .A3(new_n486_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT38), .ZN(new_n619_));
  INV_X1    g418(.A(new_n301_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n279_), .A2(new_n620_), .A3(new_n612_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT101), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n351_), .A2(new_n343_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n621_), .B2(KEYINPUT101), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n594_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n487_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n627_), .ZN(G1324gat));
  AND2_X1   g427(.A1(new_n441_), .A2(new_n495_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n617_), .A2(new_n282_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G8gat), .B1(new_n626_), .B2(new_n629_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT39), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT39), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g435(.A(new_n551_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n552_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n626_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT41), .Z(new_n642_));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n617_), .A2(new_n643_), .A3(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1326gat));
  XOR2_X1   g444(.A(new_n524_), .B(KEYINPUT102), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G22gat), .B1(new_n626_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n617_), .A2(new_n650_), .A3(new_n646_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n346_), .A2(new_n353_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n594_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT43), .B1(new_n615_), .B2(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n279_), .A2(new_n301_), .A3(new_n612_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(KEYINPUT103), .A3(KEYINPUT44), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n659_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n487_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n613_), .A2(new_n616_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n620_), .A2(new_n623_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n279_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT104), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n670_), .A2(new_n674_), .A3(new_n279_), .A4(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n303_), .A3(new_n486_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT105), .B1(new_n667_), .B2(new_n630_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n629_), .C1(new_n662_), .C2(new_n666_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n681_), .A2(new_n683_), .A3(new_n304_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n673_), .A2(new_n304_), .A3(new_n630_), .A4(new_n675_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n685_), .B(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n680_), .B1(new_n684_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n681_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n667_), .A2(KEYINPUT105), .A3(new_n630_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(G36gat), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n685_), .B(new_n688_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(G1329gat));
  OAI21_X1  g496(.A(new_n313_), .B1(new_n676_), .B2(new_n640_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n313_), .B1(new_n662_), .B2(new_n666_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n549_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(KEYINPUT109), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT109), .B1(new_n699_), .B2(new_n700_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(new_n698_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  INV_X1    g506(.A(new_n524_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G50gat), .B1(new_n668_), .B2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n677_), .A2(new_n320_), .A3(new_n646_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1331gat));
  AOI21_X1  g510(.A(new_n268_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n712_));
  NOR4_X1   g511(.A1(new_n264_), .A2(new_n266_), .A3(KEYINPUT13), .A4(new_n269_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n611_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n615_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n487_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n354_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n487_), .A2(G57gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT110), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n717_), .B2(new_n629_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT111), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n719_), .A2(G64gat), .A3(new_n629_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n717_), .B2(new_n640_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n719_), .A2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n640_), .B2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n717_), .B2(new_n647_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT112), .Z(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n719_), .A2(G78gat), .A3(new_n647_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1335gat));
  AND2_X1   g535(.A1(new_n716_), .A2(new_n671_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n486_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT113), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n715_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n301_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n486_), .A2(new_n205_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n741_), .B2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n737_), .B2(new_n630_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n629_), .A2(new_n206_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n741_), .B2(new_n745_), .ZN(G1337gat));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n221_), .A3(new_n700_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n215_), .B1(new_n741_), .B2(new_n639_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n740_), .A2(new_n301_), .A3(new_n524_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT115), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n740_), .A2(new_n756_), .A3(new_n301_), .A4(new_n524_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(G106gat), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT52), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n755_), .A2(new_n760_), .A3(G106gat), .A4(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n737_), .A2(new_n222_), .A3(new_n524_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n596_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n600_), .A2(new_n597_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n606_), .A3(new_n771_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n772_), .A2(KEYINPUT118), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(KEYINPUT118), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n608_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n248_), .A2(new_n249_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n777_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n245_), .A2(new_n255_), .A3(new_n247_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n256_), .A2(new_n778_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n263_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT56), .B(new_n263_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n611_), .A2(new_n269_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n277_), .A2(new_n775_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n769_), .B1(new_n790_), .B2(new_n624_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n787_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n778_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n250_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(new_n780_), .A3(new_n781_), .A4(new_n779_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n263_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n775_), .B(new_n270_), .C1(new_n792_), .C2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n270_), .A4(new_n775_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n655_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n773_), .A2(new_n608_), .A3(new_n774_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n612_), .A2(new_n270_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT57), .B(new_n623_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n791_), .A2(new_n801_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n301_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n611_), .B(new_n354_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(KEYINPUT116), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(KEYINPUT116), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n279_), .A2(new_n813_), .A3(new_n611_), .A4(new_n354_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(KEYINPUT54), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n811_), .A3(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n630_), .A2(new_n487_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n591_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G113gat), .B1(new_n820_), .B2(new_n612_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n823_), .A3(new_n591_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n612_), .A2(G113gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT119), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n821_), .B1(new_n825_), .B2(new_n827_), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n822_), .A2(new_n714_), .A3(new_n824_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT120), .B(G120gat), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n279_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n820_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n832_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(G1341gat));
  AOI21_X1  g634(.A(G127gat), .B1(new_n820_), .B2(new_n620_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n620_), .A2(G127gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n825_), .B2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n820_), .B2(new_n624_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n655_), .A2(G134gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n825_), .B2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n639_), .A2(new_n708_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n816_), .A2(new_n817_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT121), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n816_), .A2(new_n845_), .A3(new_n817_), .A4(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n612_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n714_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n620_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n855_));
  INV_X1    g654(.A(new_n853_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n847_), .A2(new_n620_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n855_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n847_), .B2(new_n620_), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n301_), .B(new_n853_), .C1(new_n844_), .C2(new_n846_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n847_), .B2(new_n624_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n654_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(G162gat), .B2(new_n865_), .ZN(G1347gat));
  AND2_X1   g665(.A1(new_n816_), .A2(new_n630_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n640_), .A2(new_n486_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n867_), .A2(new_n647_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n378_), .B1(new_n869_), .B2(new_n612_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n647_), .A3(new_n868_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n871_), .A2(new_n611_), .A3(new_n418_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT62), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n871_), .B2(new_n611_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1348gat));
  AOI21_X1  g676(.A(G176gat), .B1(new_n869_), .B2(new_n714_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n816_), .A2(new_n708_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n640_), .A2(new_n486_), .A3(new_n629_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n816_), .A2(KEYINPUT124), .A3(new_n708_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n279_), .A2(new_n383_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n878_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NAND4_X1  g685(.A1(new_n881_), .A2(new_n620_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n292_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n301_), .A2(new_n398_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n869_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT125), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n888_), .A2(new_n890_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1350gat));
  NAND3_X1  g694(.A1(new_n869_), .A2(new_n399_), .A3(new_n624_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G190gat), .B1(new_n871_), .B2(new_n654_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1351gat));
  NAND3_X1  g697(.A1(new_n867_), .A2(new_n487_), .A3(new_n842_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n611_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n605_), .ZN(G1352gat));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n279_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT126), .B(G204gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1353gat));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n867_), .A2(new_n487_), .A3(new_n842_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n620_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT63), .B(G211gat), .Z(new_n908_));
  NOR3_X1   g707(.A1(new_n899_), .A2(new_n301_), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT127), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n899_), .A2(new_n301_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n906_), .A2(new_n620_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n911_), .B(new_n912_), .C1(new_n913_), .C2(new_n908_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1354gat));
  AND3_X1   g714(.A1(new_n906_), .A2(G218gat), .A3(new_n655_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G218gat), .B1(new_n906_), .B2(new_n624_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


