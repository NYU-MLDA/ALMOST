//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211_));
  AOI22_X1  g010(.A1(new_n206_), .A2(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT10), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT10), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(KEYINPUT9), .A3(new_n209_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n223_), .A2(KEYINPUT68), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(KEYINPUT68), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n206_), .A2(new_n208_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT7), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n227_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n230_), .A2(new_n216_), .A3(new_n213_), .A4(KEYINPUT64), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n221_), .A2(new_n209_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n236_));
  OAI22_X1  g035(.A1(new_n224_), .A2(new_n225_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT15), .ZN(new_n238_));
  OR2_X1    g037(.A1(G29gat), .A2(G36gat), .ZN(new_n239_));
  INV_X1    g038(.A(G43gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G29gat), .A2(G36gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G50gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n240_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G43gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(G50gat), .B1(new_n248_), .B2(new_n242_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n238_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(G50gat), .A3(new_n242_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT15), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n204_), .B1(new_n237_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n246_), .A2(new_n249_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n256_), .B(new_n223_), .C1(new_n236_), .C2(new_n235_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n236_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n262_), .A2(KEYINPUT72), .A3(new_n256_), .A4(new_n223_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n255_), .A2(KEYINPUT74), .A3(new_n259_), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT71), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n255_), .A2(KEYINPUT73), .A3(new_n259_), .A4(new_n263_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT75), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G134gat), .ZN(new_n276_));
  INV_X1    g075(.A(G162gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT36), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n270_), .A2(new_n280_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n274_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n278_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT36), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n270_), .A2(new_n284_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT37), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n279_), .ZN(new_n290_));
  OAI211_X1 g089(.A(KEYINPUT37), .B(new_n285_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G127gat), .B(G155gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G183gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G211gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT67), .B1(new_n297_), .B2(KEYINPUT17), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n298_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G71gat), .ZN(new_n309_));
  INV_X1    g108(.A(G78gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G71gat), .A2(G78gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G57gat), .B(G64gat), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(new_n312_), .C1(new_n313_), .C2(KEYINPUT11), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT66), .ZN(new_n315_));
  AND2_X1   g114(.A1(G57gat), .A2(G64gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G57gat), .A2(G64gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n311_), .A4(new_n312_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n318_), .A2(new_n319_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n315_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n315_), .B2(new_n322_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n298_), .A2(new_n307_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n308_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n308_), .B2(new_n327_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n293_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT76), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(KEYINPUT85), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(new_n343_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n338_), .B(new_n339_), .C1(new_n342_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n340_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n336_), .B(KEYINPUT84), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n339_), .B(KEYINPUT1), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n349_), .B(new_n344_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G120gat), .ZN(new_n354_));
  AND2_X1   g153(.A1(G127gat), .A2(G134gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G127gat), .A2(G134gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT82), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G127gat), .ZN(new_n358_));
  INV_X1    g157(.A(G134gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G127gat), .A2(G134gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G113gat), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n357_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n357_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n354_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n355_), .A2(new_n356_), .A3(KEYINPUT82), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n361_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n369_));
  OAI21_X1  g168(.A(G113gat), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n357_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(G120gat), .A3(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n367_), .A2(KEYINPUT83), .A3(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT83), .B1(new_n367_), .B2(new_n372_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n335_), .B(new_n353_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT97), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT96), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n367_), .A2(new_n372_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n353_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n367_), .A2(new_n372_), .A3(KEYINPUT83), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n381_), .B1(new_n385_), .B2(new_n353_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n379_), .B1(new_n386_), .B2(KEYINPUT4), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n383_), .A2(new_n384_), .B1(new_n352_), .B2(new_n348_), .ZN(new_n388_));
  NOR4_X1   g187(.A1(new_n388_), .A2(new_n381_), .A3(KEYINPUT95), .A4(new_n335_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n376_), .B(new_n378_), .C1(new_n387_), .C2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n378_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT98), .B(G85gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT0), .B(G57gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n396_), .B(new_n397_), .Z(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n390_), .A2(new_n392_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(KEYINPUT100), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n390_), .A2(new_n403_), .A3(new_n392_), .A4(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  OR2_X1    g205(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT77), .B(G183gat), .Z(new_n408_));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G190gat), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(KEYINPUT26), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(KEYINPUT26), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT78), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G169gat), .ZN(new_n416_));
  INV_X1    g215(.A(G176gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT24), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G169gat), .A2(G176gat), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n421_), .A2(KEYINPUT79), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT80), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G183gat), .A3(G190gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(KEYINPUT23), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT79), .B1(new_n421_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n415_), .A2(new_n422_), .A3(new_n430_), .A4(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n427_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n423_), .A2(KEYINPUT23), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT81), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n435_), .A2(KEYINPUT81), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n436_), .A2(new_n437_), .B1(new_n411_), .B2(new_n408_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G169gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n433_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G197gat), .A2(G204gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT87), .B(G197gat), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT21), .B(new_n443_), .C1(new_n444_), .C2(G204gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(G211gat), .B(G218gat), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G204gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G197gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n445_), .B(new_n447_), .C1(new_n450_), .C2(KEYINPUT21), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(KEYINPUT21), .A3(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n406_), .B1(new_n442_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT25), .B(G183gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT91), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n412_), .A2(new_n413_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n456_), .A2(new_n457_), .B1(new_n420_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n436_), .A2(new_n437_), .ZN(new_n460_));
  OR3_X1    g259(.A1(new_n458_), .A2(new_n420_), .A3(new_n418_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n453_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n430_), .B1(G183gat), .B2(G190gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n440_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n454_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT19), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n442_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n463_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n462_), .A2(new_n465_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n453_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n473_), .A2(KEYINPUT20), .A3(new_n469_), .A4(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484_));
  INV_X1    g283(.A(new_n482_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n471_), .A2(new_n476_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(KEYINPUT94), .A3(new_n482_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(new_n469_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n473_), .A2(KEYINPUT20), .A3(new_n475_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n469_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n485_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(KEYINPUT27), .A3(new_n483_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT31), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n442_), .A2(new_n384_), .A3(new_n383_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n442_), .B1(new_n384_), .B2(new_n383_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n498_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n472_), .A2(new_n385_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n498_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G99gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT30), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(new_n510_), .A3(new_n505_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n515_));
  XOR2_X1   g314(.A(G22gat), .B(G50gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n515_), .B(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G78gat), .B(G106gat), .Z(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT88), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n463_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n521_), .B(KEYINPUT88), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n453_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n520_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n519_), .B1(new_n530_), .B2(KEYINPUT89), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT90), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n525_), .A2(new_n529_), .A3(new_n520_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n530_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n535_), .B(new_n519_), .C1(new_n530_), .C2(KEYINPUT89), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n514_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n512_), .A2(new_n513_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n537_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n538_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n405_), .A2(new_n496_), .A3(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(new_n538_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n493_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n493_), .A2(KEYINPUT99), .A3(new_n548_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n402_), .A2(new_n404_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT33), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n401_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n487_), .A2(new_n488_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n376_), .B(new_n391_), .C1(new_n387_), .C2(new_n389_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n386_), .A2(new_n378_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n398_), .A3(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n390_), .A2(KEYINPUT33), .A3(new_n392_), .A4(new_n400_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n556_), .A2(new_n557_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n546_), .B1(new_n554_), .B2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n545_), .B1(new_n563_), .B2(new_n514_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n256_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(new_n305_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n254_), .A2(new_n305_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n256_), .B(new_n305_), .Z(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(G229gat), .A3(G233gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n416_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(G197gat), .Z(new_n576_));
  OR2_X1    g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n576_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n581_));
  INV_X1    g380(.A(G230gat), .ZN(new_n582_));
  INV_X1    g381(.A(G233gat), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT67), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n315_), .A2(new_n322_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n323_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n315_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(KEYINPUT67), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n223_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n586_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n584_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n237_), .B(KEYINPUT12), .C1(new_n324_), .C2(new_n325_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n594_), .B(new_n598_), .C1(new_n596_), .C2(KEYINPUT12), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n599_), .B2(new_n584_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n597_), .B(new_n607_), .C1(new_n599_), .C2(new_n584_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n606_), .A2(KEYINPUT13), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT13), .B1(new_n606_), .B2(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n581_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n596_), .A2(KEYINPUT12), .ZN(new_n614_));
  INV_X1    g413(.A(new_n584_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n594_), .A4(new_n598_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n607_), .B1(new_n616_), .B2(new_n597_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n608_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n613_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n606_), .A2(KEYINPUT13), .A3(new_n608_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT70), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n612_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n564_), .A2(new_n580_), .A3(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n334_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n405_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n300_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  INV_X1    g428(.A(new_n286_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n331_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n625_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(new_n627_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n300_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n496_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n301_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT39), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n626_), .A2(new_n301_), .A3(new_n635_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n626_), .A2(new_n642_), .A3(new_n541_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT102), .Z(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n632_), .B2(new_n541_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1326gat));
  INV_X1    g446(.A(G22gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n632_), .B2(new_n546_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT42), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n626_), .A2(new_n648_), .A3(new_n546_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1327gat));
  NOR2_X1   g451(.A1(new_n624_), .A2(new_n580_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n331_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT103), .B(KEYINPUT43), .C1(new_n564_), .C2(new_n293_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n541_), .B(new_n546_), .C1(new_n554_), .C2(new_n562_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n292_), .B1(new_n658_), .B2(new_n545_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT43), .B1(new_n659_), .B2(KEYINPUT103), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n554_), .A2(new_n562_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n546_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n514_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n545_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n293_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n656_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n663_), .A2(new_n627_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n663_), .A2(KEYINPUT104), .A3(new_n627_), .A4(new_n673_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(G29gat), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n630_), .A2(new_n331_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT105), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n625_), .A2(new_n680_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n681_), .A2(G29gat), .A3(new_n405_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n678_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(KEYINPUT106), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1328gat));
  NOR3_X1   g486(.A1(new_n681_), .A2(G36gat), .A3(new_n496_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT45), .Z(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n663_), .A2(new_n635_), .A3(new_n673_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n689_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(G1329gat));
  OAI21_X1  g495(.A(new_n240_), .B1(new_n681_), .B2(new_n514_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT109), .Z(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n655_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n662_), .B(new_n654_), .C1(new_n671_), .C2(new_n656_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n240_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT108), .B1(new_n701_), .B2(new_n541_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n663_), .A2(G43gat), .A3(new_n541_), .A4(new_n673_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n702_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT47), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n708_), .B(new_n698_), .C1(new_n702_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n663_), .A2(new_n546_), .A3(new_n673_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n663_), .A2(new_n713_), .A3(new_n546_), .A4(new_n673_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(G50gat), .A3(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n625_), .A2(new_n244_), .A3(new_n546_), .A4(new_n680_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n719_), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1331gat));
  NOR2_X1   g520(.A1(new_n623_), .A2(new_n579_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n564_), .A2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n334_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n627_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n724_), .A2(new_n631_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n627_), .A2(G57gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  INV_X1    g528(.A(G64gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n730_), .A3(new_n635_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n635_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G64gat), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT48), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT48), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n725_), .A2(new_n309_), .A3(new_n541_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n727_), .A2(new_n541_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G71gat), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT49), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT49), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1334gat));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n310_), .A3(new_n546_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n727_), .A2(new_n546_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G78gat), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT50), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(KEYINPUT50), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n724_), .A2(new_n680_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n627_), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n332_), .B(new_n723_), .C1(new_n671_), .C2(new_n656_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n405_), .A2(new_n219_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  OAI21_X1  g553(.A(new_n220_), .B1(new_n749_), .B2(new_n496_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT112), .ZN(new_n756_));
  INV_X1    g555(.A(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n635_), .A2(G92gat), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT113), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT114), .ZN(G1337gat));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n752_), .A2(new_n541_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G99gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n541_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n749_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n762_), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT115), .B(new_n766_), .C1(new_n763_), .C2(G99gat), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n768_), .A2(new_n770_), .A3(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n750_), .A2(new_n213_), .A3(new_n546_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n752_), .A2(new_n546_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(G106gat), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT52), .B(new_n213_), .C1(new_n752_), .C2(new_n546_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n609_), .A2(new_n610_), .A3(new_n579_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n288_), .A2(new_n332_), .A3(new_n291_), .A4(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  NOR2_X1   g587(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n788_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n785_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT37), .B1(new_n282_), .B2(new_n285_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n619_), .A2(new_n580_), .A3(new_n620_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n291_), .ZN(new_n796_));
  NOR4_X1   g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .A4(new_n331_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT117), .B1(new_n797_), .B2(new_n789_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n785_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n793_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n571_), .A2(new_n569_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n568_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n576_), .B(new_n804_), .C1(new_n805_), .C2(new_n569_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n577_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n599_), .A2(new_n584_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT55), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n616_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n599_), .A2(new_n813_), .A3(new_n584_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n605_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n599_), .B2(new_n584_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n599_), .A2(new_n584_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT56), .B(new_n605_), .C1(new_n820_), .C2(new_n814_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n817_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n579_), .A2(new_n608_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n809_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n286_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n605_), .B1(new_n820_), .B2(new_n814_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n829_), .B2(new_n821_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT57), .B(new_n286_), .C1(new_n830_), .C2(new_n808_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n826_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n807_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n608_), .B(new_n835_), .C1(new_n817_), .C2(new_n822_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n829_), .A2(new_n821_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n608_), .A4(new_n835_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n292_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n286_), .B1(new_n830_), .B2(new_n808_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n331_), .B1(new_n834_), .B2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n802_), .A2(new_n803_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n803_), .B1(new_n802_), .B2(new_n846_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n635_), .A2(new_n405_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n543_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n847_), .A2(new_n848_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853_), .B2(new_n579_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n802_), .A2(new_n846_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n851_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT121), .B(new_n858_), .C1(new_n853_), .C2(new_n859_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n580_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n854_), .B1(new_n864_), .B2(G113gat), .ZN(G1340gat));
  XNOR2_X1  g664(.A(KEYINPUT122), .B(G120gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n860_), .B2(new_n623_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n624_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n853_), .B(new_n870_), .C1(new_n869_), .C2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n867_), .A2(new_n873_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n853_), .B2(new_n332_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n331_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n853_), .B2(new_n630_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n293_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n847_), .A2(new_n848_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n540_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n849_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n579_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n624_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g687(.A1(new_n883_), .A2(new_n331_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT61), .B(G155gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT124), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n889_), .B(new_n891_), .ZN(G1346gat));
  NOR3_X1   g691(.A1(new_n883_), .A2(new_n277_), .A3(new_n293_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n884_), .A2(new_n630_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n277_), .B2(new_n894_), .ZN(G1347gat));
  INV_X1    g694(.A(new_n855_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n635_), .A2(new_n405_), .A3(new_n541_), .A4(new_n666_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n579_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899_), .B2(KEYINPUT62), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT62), .B1(new_n899_), .B2(KEYINPUT22), .ZN(new_n901_));
  MUX2_X1   g700(.A(G169gat), .B(new_n900_), .S(new_n901_), .Z(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n898_), .B2(new_n624_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n847_), .A2(new_n848_), .A3(new_n897_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n623_), .A2(new_n417_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  INV_X1    g705(.A(new_n898_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n907_), .A2(new_n456_), .A3(new_n331_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n332_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n408_), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n907_), .B2(new_n293_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n898_), .A2(new_n457_), .A3(new_n630_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1351gat));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n405_), .A2(new_n882_), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n915_), .B(KEYINPUT125), .Z(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n496_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n881_), .A2(new_n914_), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n855_), .A2(KEYINPUT119), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n802_), .A2(new_n846_), .A3(new_n803_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n579_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n624_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g726(.A(KEYINPUT63), .B(G211gat), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n914_), .B1(new_n881_), .B2(new_n917_), .ZN(new_n929_));
  AND4_X1   g728(.A1(new_n914_), .A2(new_n919_), .A3(new_n920_), .A4(new_n917_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n332_), .B(new_n928_), .C1(new_n929_), .C2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n332_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n923_), .A2(KEYINPUT127), .A3(new_n332_), .A4(new_n928_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n933_), .A2(new_n936_), .A3(new_n937_), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n923_), .B2(new_n630_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n293_), .B1(new_n918_), .B2(new_n922_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(G218gat), .B2(new_n940_), .ZN(G1355gat));
endmodule


