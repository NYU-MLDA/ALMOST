//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(new_n203_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT91), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n208_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n211_), .B(new_n214_), .C1(new_n209_), .C2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT92), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n203_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n204_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(new_n206_), .B2(new_n223_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(G183gat), .B2(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n216_), .A3(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  INV_X1    g028(.A(G218gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(G211gat), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G197gat), .B(G204gat), .Z(new_n232_));
  OAI221_X1 g031(.A(new_n231_), .B1(G211gat), .B2(new_n230_), .C1(new_n232_), .C2(KEYINPUT21), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n202_), .B1(new_n228_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G226gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT19), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n235_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G169gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n207_), .B2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n214_), .A2(new_n245_), .ZN(new_n246_));
  OAI221_X1 g045(.A(new_n225_), .B1(KEYINPUT24), .B2(new_n215_), .C1(new_n246_), .C2(KEYINPUT83), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(KEYINPUT83), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n240_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT93), .Z(new_n251_));
  NAND3_X1  g050(.A1(new_n236_), .A2(new_n239_), .A3(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n228_), .A2(new_n235_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT20), .B1(new_n240_), .B2(new_n249_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n238_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G64gat), .B(G92gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT27), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT97), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n239_), .B1(new_n236_), .B2(new_n251_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n253_), .A2(new_n238_), .A3(new_n254_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n260_), .B(KEYINPUT96), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n265_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  OAI211_X1 g070(.A(KEYINPUT97), .B(new_n271_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n263_), .A2(KEYINPUT27), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n264_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n276_), .A2(KEYINPUT86), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(KEYINPUT86), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G113gat), .B(G120gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G155gat), .ZN(new_n285_));
  INV_X1    g084(.A(G162gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n285_), .A2(new_n286_), .A3(KEYINPUT1), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(KEYINPUT3), .ZN(new_n293_));
  OR3_X1    g092(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n298_), .B(new_n284_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n292_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n281_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT4), .ZN(new_n302_));
  INV_X1    g101(.A(new_n300_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n281_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT94), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G29gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G85gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G57gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n281_), .B(KEYINPUT31), .Z(new_n320_));
  XOR2_X1   g119(.A(new_n249_), .B(KEYINPUT30), .Z(new_n321_));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G43gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(G15gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n325_), .B(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n323_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n322_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n321_), .A2(new_n322_), .A3(new_n329_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n320_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n320_), .A3(new_n333_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n235_), .B1(new_n303_), .B2(KEYINPUT29), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n300_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT28), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n300_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT89), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n347_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n340_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n339_), .B(KEYINPUT89), .C1(new_n348_), .C2(new_n349_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G78gat), .B(G106gat), .Z(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n335_), .B(new_n336_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n359_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n336_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n357_), .C1(new_n363_), .C2(new_n334_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n275_), .B(new_n319_), .C1(new_n361_), .C2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n302_), .A2(new_n306_), .A3(new_n305_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n301_), .A2(new_n307_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n315_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT33), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n308_), .A2(KEYINPUT33), .A3(new_n309_), .A4(new_n314_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n370_), .A2(new_n317_), .B1(new_n371_), .B2(KEYINPUT95), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n371_), .A2(KEYINPUT95), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n262_), .A3(new_n263_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n252_), .A2(new_n255_), .A3(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(new_n318_), .C1(new_n268_), .C2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n358_), .A2(new_n359_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n363_), .A2(new_n334_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n366_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G1gat), .ZN(new_n383_));
  INV_X1    g182(.A(G8gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT14), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT79), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(KEYINPUT79), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G15gat), .B(G22gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G1gat), .B(G8gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT80), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n389_), .B(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G29gat), .B(G36gat), .Z(new_n393_));
  XOR2_X1   g192(.A(G43gat), .B(G50gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n395_), .B(KEYINPUT15), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G229gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT82), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n392_), .B(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n402_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n397_), .A2(new_n399_), .A3(new_n406_), .A4(new_n401_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G113gat), .B(G141gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G169gat), .B(G197gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT98), .B1(new_n382_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n417_));
  INV_X1    g216(.A(new_n415_), .ZN(new_n418_));
  AOI211_X1 g217(.A(new_n417_), .B(new_n418_), .C1(new_n366_), .C2(new_n381_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n421_));
  NAND2_X1  g220(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G85gat), .B(G92gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT6), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(G99gat), .A3(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  AOI211_X1 g232(.A(new_n423_), .B(new_n424_), .C1(new_n428_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT7), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n431_), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n429_), .A2(KEYINPUT6), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n425_), .B(new_n438_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n424_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n422_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT71), .B1(new_n434_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n430_), .A2(new_n432_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n425_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n423_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n422_), .A3(new_n442_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n444_), .A2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n455_), .A2(new_n437_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT65), .B(G85gat), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT66), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G92gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n457_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT9), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(G85gat), .B2(G92gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n456_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT72), .B1(new_n452_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT72), .ZN(new_n470_));
  INV_X1    g269(.A(new_n468_), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n470_), .B(new_n471_), .C1(new_n444_), .C2(new_n451_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n398_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT74), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n468_), .B1(new_n434_), .B2(new_n443_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT68), .B(new_n468_), .C1(new_n434_), .C2(new_n443_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n395_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n473_), .A2(new_n474_), .A3(new_n480_), .A4(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n473_), .A2(new_n474_), .A3(new_n480_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n483_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT35), .B1(new_n473_), .B2(new_n480_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G190gat), .B(G218gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT75), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G134gat), .B(G162gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT36), .Z(new_n494_));
  AOI21_X1  g293(.A(new_n421_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n493_), .A2(KEYINPUT36), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n485_), .B(new_n497_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n489_), .A2(new_n421_), .A3(new_n494_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n494_), .B(KEYINPUT76), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n489_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n498_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT37), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n508_), .B1(new_n479_), .B2(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT69), .B(new_n515_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n477_), .A2(new_n515_), .A3(new_n478_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT70), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n507_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(KEYINPUT12), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n507_), .B1(new_n479_), .B2(new_n516_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n521_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n528_), .B1(new_n521_), .B2(new_n529_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n526_), .B(new_n527_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n523_), .A2(new_n532_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT13), .B1(new_n538_), .B2(new_n540_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n515_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n392_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT16), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n552_), .B(KEYINPUT17), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n548_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n506_), .A2(new_n545_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT81), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(KEYINPUT81), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n319_), .A2(G1gat), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n420_), .A2(new_n561_), .A3(new_n562_), .A4(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT38), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT99), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n499_), .A2(new_n498_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(new_n495_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n366_), .B2(new_n381_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n545_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n571_), .A2(new_n558_), .A3(new_n418_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT100), .Z(new_n574_));
  AOI21_X1  g373(.A(new_n383_), .B1(new_n574_), .B2(new_n318_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT101), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n564_), .A2(new_n565_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT102), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n567_), .A2(new_n577_), .A3(new_n579_), .ZN(G1324gat));
  AND3_X1   g379(.A1(new_n420_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n275_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n384_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n573_), .A2(KEYINPUT103), .A3(new_n275_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n585_), .A2(G8gat), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT103), .B1(new_n573_), .B2(new_n275_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n584_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AND4_X1   g387(.A1(new_n584_), .A2(new_n585_), .A3(G8gat), .A4(new_n587_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n583_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT40), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n583_), .B(KEYINPUT40), .C1(new_n588_), .C2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1325gat));
  INV_X1    g393(.A(new_n380_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n327_), .B1(new_n574_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n581_), .A2(new_n327_), .A3(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1326gat));
  INV_X1    g399(.A(G22gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n379_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n574_), .B2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT42), .Z(new_n604_));
  NAND3_X1  g403(.A1(new_n581_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1327gat));
  INV_X1    g405(.A(new_n569_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n571_), .A2(new_n559_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT107), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT107), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n611_), .B(new_n608_), .C1(new_n416_), .C2(new_n419_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(G29gat), .B1(new_n613_), .B2(new_n318_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n571_), .A2(new_n559_), .A3(new_n418_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n506_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n382_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT43), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  AOI211_X1 g419(.A(KEYINPUT105), .B(new_n620_), .C1(new_n382_), .C2(new_n616_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT44), .B(new_n615_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n615_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n620_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT43), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n622_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n318_), .A2(G29gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n614_), .B1(new_n630_), .B2(new_n631_), .ZN(G1328gat));
  NOR2_X1   g431(.A1(new_n275_), .A2(G36gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n610_), .A2(new_n612_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT45), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT45), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n610_), .A2(new_n636_), .A3(new_n612_), .A4(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n622_), .B(new_n582_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G36gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n638_), .B(new_n640_), .C1(KEYINPUT108), .C2(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1329gat));
  NAND3_X1  g444(.A1(new_n610_), .A2(new_n595_), .A3(new_n612_), .ZN(new_n646_));
  INV_X1    g445(.A(G43gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n595_), .A2(G43gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n629_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g450(.A(G50gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n613_), .A2(new_n652_), .A3(new_n602_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n622_), .B(new_n602_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT109), .B1(new_n654_), .B2(G50gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1331gat));
  NAND2_X1  g456(.A1(new_n571_), .A2(new_n418_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n366_), .B2(new_n381_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n659_), .A2(new_n559_), .A3(new_n506_), .ZN(new_n660_));
  INV_X1    g459(.A(G57gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n318_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n570_), .A2(new_n559_), .A3(new_n571_), .A4(new_n418_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n319_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1332gat));
  OAI21_X1  g464(.A(G64gat), .B1(new_n663_), .B2(new_n275_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT48), .ZN(new_n667_));
  INV_X1    g466(.A(G64gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n668_), .A3(new_n582_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n663_), .B2(new_n380_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G71gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n674_), .A3(new_n595_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1334gat));
  OAI21_X1  g475(.A(G78gat), .B1(new_n663_), .B2(new_n379_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT50), .ZN(new_n678_));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n660_), .A2(new_n679_), .A3(new_n602_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1335gat));
  AND3_X1   g480(.A1(new_n659_), .A2(new_n558_), .A3(new_n569_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G85gat), .B1(new_n682_), .B2(new_n318_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n625_), .A2(new_n626_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n658_), .A2(new_n559_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n318_), .A2(new_n458_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n683_), .B1(new_n687_), .B2(new_n688_), .ZN(G1336gat));
  AOI21_X1  g488(.A(G92gat), .B1(new_n682_), .B2(new_n582_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n275_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n687_), .B2(new_n691_), .ZN(G1337gat));
  OAI21_X1  g491(.A(G99gat), .B1(new_n686_), .B2(new_n380_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n380_), .A2(new_n454_), .A3(new_n453_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n682_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(KEYINPUT111), .A3(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g496(.A1(new_n682_), .A2(new_n437_), .A3(new_n602_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n602_), .B(new_n685_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT52), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(G106gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G106gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g503(.A1(new_n582_), .A2(new_n319_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n365_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n532_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT55), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT55), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n532_), .A2(new_n707_), .A3(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n519_), .B(new_n526_), .C1(new_n531_), .C2(new_n530_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n507_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n711_), .A3(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT114), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT114), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n714_), .A2(new_n717_), .A3(KEYINPUT56), .A4(new_n537_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n537_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT56), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n718_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n411_), .B1(new_n404_), .B2(new_n401_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n401_), .B2(new_n400_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n414_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT113), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n540_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n722_), .A2(KEYINPUT58), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT58), .B1(new_n722_), .B2(new_n727_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n506_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n540_), .A2(new_n415_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n721_), .B2(new_n715_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n541_), .A2(new_n726_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n607_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n732_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n708_), .A2(KEYINPUT55), .B1(new_n712_), .B2(new_n507_), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n720_), .B(new_n539_), .C1(new_n740_), .C2(new_n711_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n537_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n734_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT57), .A3(new_n607_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n738_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n558_), .B1(new_n731_), .B2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n506_), .A2(new_n545_), .A3(new_n559_), .A4(new_n418_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT54), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n706_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G113gat), .B1(new_n750_), .B2(new_n415_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n749_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n706_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT59), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT59), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT115), .B1(new_n750_), .B2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT57), .B1(new_n744_), .B2(new_n607_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n737_), .B(new_n569_), .C1(new_n743_), .C2(new_n734_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n722_), .A2(new_n727_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n616_), .A3(new_n728_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n559_), .B1(new_n760_), .B2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n748_), .B(KEYINPUT54), .Z(new_n766_));
  OAI211_X1 g565(.A(new_n756_), .B(new_n753_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n755_), .B1(new_n757_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n750_), .A2(KEYINPUT115), .A3(new_n756_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n767_), .A2(new_n768_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT116), .A3(new_n755_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n415_), .A2(G113gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT117), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n751_), .B1(new_n777_), .B2(new_n779_), .ZN(G1340gat));
  INV_X1    g579(.A(G120gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n571_), .B1(new_n750_), .B2(new_n756_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n775_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n781_), .A2(KEYINPUT60), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT60), .ZN(new_n786_));
  AOI21_X1  g585(.A(G120gat), .B1(new_n571_), .B2(new_n786_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n754_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT118), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790_));
  INV_X1    g589(.A(new_n788_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n782_), .B1(new_n774_), .B2(new_n773_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n790_), .B(new_n791_), .C1(new_n792_), .C2(new_n781_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(G1341gat));
  AOI21_X1  g593(.A(G127gat), .B1(new_n750_), .B2(new_n559_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT119), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n559_), .A2(G127gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n777_), .B2(new_n797_), .ZN(G1342gat));
  AOI21_X1  g597(.A(G134gat), .B1(new_n750_), .B2(new_n569_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n616_), .A2(G134gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n777_), .B2(new_n800_), .ZN(G1343gat));
  NAND3_X1  g600(.A1(new_n752_), .A2(new_n361_), .A3(new_n705_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n418_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n545_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT120), .B(G148gat), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1345gat));
  NOR2_X1   g606(.A1(new_n802_), .A2(new_n558_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  NOR3_X1   g609(.A1(new_n802_), .A2(new_n286_), .A3(new_n506_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n802_), .A2(new_n607_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(G162gat), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n813_), .A2(KEYINPUT121), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(KEYINPUT121), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(G1347gat));
  AOI21_X1  g615(.A(new_n602_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n275_), .A2(new_n318_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n595_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT122), .B1(new_n821_), .B2(new_n418_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n817_), .A2(new_n823_), .A3(new_n415_), .A4(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(G169gat), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n817_), .A2(new_n820_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n415_), .A3(new_n220_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n822_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n824_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n829_), .A3(new_n830_), .ZN(G1348gat));
  AOI21_X1  g630(.A(G176gat), .B1(new_n828_), .B2(new_n571_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n817_), .B(KEYINPUT123), .Z(new_n833_));
  NOR3_X1   g632(.A1(new_n819_), .A2(new_n221_), .A3(new_n545_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(G1349gat));
  NOR3_X1   g634(.A1(new_n821_), .A2(new_n558_), .A3(new_n212_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n559_), .A3(new_n820_), .ZN(new_n837_));
  INV_X1    g636(.A(G183gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1350gat));
  NAND3_X1  g638(.A1(new_n828_), .A2(new_n569_), .A3(new_n213_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G190gat), .B1(new_n821_), .B2(new_n506_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT124), .ZN(G1351gat));
  NAND3_X1  g642(.A1(new_n752_), .A2(new_n361_), .A3(new_n818_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n752_), .A2(KEYINPUT125), .A3(new_n361_), .A4(new_n818_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n415_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n571_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g651(.A(new_n558_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT126), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n854_), .B(new_n856_), .ZN(G1354gat));
  AOI211_X1 g656(.A(new_n230_), .B(new_n506_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n607_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT127), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G218gat), .B1(new_n859_), .B2(new_n860_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n858_), .B1(new_n861_), .B2(new_n862_), .ZN(G1355gat));
endmodule


