//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT76), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT76), .B1(new_n204_), .B2(new_n206_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(G134gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n203_), .A2(G127gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT76), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n216_), .A3(KEYINPUT77), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n218_), .B(new_n202_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n220_), .B(KEYINPUT78), .Z(new_n221_));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n224_), .A2(G169gat), .B1(new_n225_), .B2(new_n222_), .ZN(new_n226_));
  OR2_X1    g025(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n226_), .B1(new_n230_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT25), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n229_), .A2(KEYINPUT26), .ZN(new_n242_));
  NOR2_X1   g041(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n241_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n233_), .A2(new_n234_), .ZN(new_n246_));
  INV_X1    g045(.A(G169gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n223_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT24), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n225_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n236_), .B1(new_n245_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G71gat), .B(G99gat), .ZN(new_n255_));
  INV_X1    g054(.A(G43gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n254_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n221_), .B(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(G15gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT30), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT31), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n259_), .B(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G141gat), .B(G148gat), .Z(new_n266_));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n267_), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT80), .B1(new_n267_), .B2(KEYINPUT1), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n271_));
  INV_X1    g070(.A(G155gat), .ZN(new_n272_));
  INV_X1    g071(.A(G162gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G155gat), .A3(G162gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n266_), .B1(new_n270_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT81), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT3), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n287_), .A2(new_n283_), .A3(new_n284_), .A4(KEYINPUT81), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n274_), .A2(new_n267_), .A3(new_n277_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n279_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT28), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n279_), .A2(new_n291_), .A3(new_n295_), .A4(new_n292_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G22gat), .B(G50gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G228gat), .A2(G233gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n292_), .B1(new_n279_), .B2(new_n291_), .ZN(new_n303_));
  OR2_X1    g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT21), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(KEYINPUT21), .A3(new_n305_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n302_), .B1(new_n303_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n267_), .A2(KEYINPUT1), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n267_), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n322_), .A2(new_n266_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n301_), .B(new_n313_), .C1(new_n323_), .C2(new_n292_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT82), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT83), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n315_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT84), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n315_), .A2(new_n324_), .A3(new_n330_), .A4(new_n327_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n315_), .A2(new_n324_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n326_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n300_), .A2(new_n329_), .A3(new_n331_), .A4(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n328_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n336_));
  OAI22_X1  g135(.A1(new_n335_), .A2(new_n336_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G85gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT0), .B(G57gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n279_), .A2(new_n291_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n220_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n209_), .A2(new_n216_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n323_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n217_), .A2(new_n219_), .B1(new_n279_), .B2(new_n291_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n345_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n343_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n346_), .A2(new_n279_), .A3(new_n291_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n350_), .A2(new_n359_), .A3(new_n351_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n220_), .A2(new_n351_), .A3(new_n344_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n349_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT89), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n343_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n355_), .A4(new_n354_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n265_), .A2(new_n339_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n371_));
  AND2_X1   g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  AOI211_X1 g172(.A(new_n370_), .B(new_n373_), .C1(new_n254_), .C2(new_n313_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n251_), .A2(KEYINPUT86), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT24), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n225_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n248_), .A2(new_n375_), .A3(new_n377_), .A4(new_n249_), .ZN(new_n380_));
  AND2_X1   g179(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n238_), .B(new_n240_), .C1(new_n381_), .C2(new_n243_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n379_), .A2(new_n246_), .A3(new_n380_), .A4(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n247_), .A2(KEYINPUT22), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n222_), .A2(G169gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT87), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT87), .B1(new_n385_), .B2(new_n386_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n223_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n233_), .B(new_n234_), .C1(G183gat), .C2(G190gat), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n391_), .A2(new_n249_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n384_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT87), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n222_), .A2(G169gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n247_), .A2(KEYINPUT22), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(G176gat), .B1(new_n397_), .B2(new_n387_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(new_n249_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n398_), .A2(new_n399_), .A3(KEYINPUT88), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n314_), .B(new_n383_), .C1(new_n393_), .C2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n374_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT20), .B1(new_n254_), .B2(new_n313_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n383_), .B1(new_n393_), .B2(new_n400_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n313_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n373_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n402_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT18), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n246_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n241_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT26), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n416_), .B1(new_n418_), .B2(new_n243_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n246_), .B1(G183gat), .B2(new_n229_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n415_), .A2(new_n419_), .B1(new_n420_), .B2(new_n226_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n370_), .B1(new_n421_), .B2(new_n314_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n383_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n390_), .A2(new_n392_), .A3(new_n384_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT88), .B1(new_n398_), .B2(new_n399_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n422_), .B1(new_n426_), .B2(new_n314_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n427_), .A2(new_n373_), .B1(new_n401_), .B2(new_n374_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n413_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n414_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n413_), .B(KEYINPUT95), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n383_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT92), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n383_), .B(new_n437_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n314_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n370_), .B1(new_n254_), .B2(new_n313_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n406_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n441_), .A2(new_n442_), .B1(new_n427_), .B2(new_n373_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT93), .B(new_n406_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n434_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n445_), .A2(KEYINPUT96), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT96), .B1(new_n445_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n433_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT99), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(KEYINPUT99), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n369_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n338_), .A2(new_n366_), .A3(new_n358_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n433_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT98), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n445_), .A2(new_n447_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n445_), .A2(KEYINPUT96), .A3(new_n447_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT98), .A3(new_n454_), .A4(new_n433_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n366_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n343_), .A2(new_n465_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n364_), .A2(new_n355_), .A3(new_n354_), .A4(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n348_), .A2(new_n349_), .A3(new_n361_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n345_), .A2(new_n347_), .A3(new_n362_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n343_), .A3(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n414_), .A3(new_n430_), .A4(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT90), .B1(new_n467_), .B2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n414_), .A2(new_n430_), .A3(new_n472_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n466_), .A4(new_n469_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT32), .B(new_n429_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT91), .B1(new_n413_), .B2(new_n479_), .ZN(new_n480_));
  OR3_X1    g279(.A1(new_n413_), .A2(KEYINPUT91), .A3(new_n479_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n428_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n367_), .A2(new_n478_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n339_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT94), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n487_), .A3(new_n339_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n464_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n265_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n453_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G29gat), .B(G36gat), .Z(new_n492_));
  XOR2_X1   g291(.A(G43gat), .B(G50gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G8gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  OR2_X1    g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n494_), .B(KEYINPUT73), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n503_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n505_), .B(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(new_n507_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G113gat), .B(G141gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT74), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G169gat), .B(G197gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n511_), .B(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n491_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT6), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(G99gat), .A3(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G85gat), .B(G92gat), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT64), .B(G92gat), .Z(new_n531_));
  INV_X1    g330(.A(KEYINPUT9), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(G85gat), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n525_), .A2(new_n528_), .A3(new_n530_), .A4(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT7), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n525_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n523_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n535_), .B1(new_n540_), .B2(new_n529_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n534_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G78gat), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n542_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n549_), .B(new_n534_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n518_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT12), .B1(new_n542_), .B2(new_n550_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n534_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n539_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT66), .ZN(new_n559_));
  INV_X1    g358(.A(new_n541_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT66), .B1(new_n539_), .B2(new_n541_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n550_), .A2(KEYINPUT12), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n556_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n552_), .A2(new_n566_), .A3(new_n518_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n552_), .B2(new_n518_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n554_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n575_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n577_), .A2(KEYINPUT68), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT68), .B1(new_n577_), .B2(new_n578_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G190gat), .B(G218gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT71), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n563_), .A2(new_n496_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT70), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT35), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n494_), .B(new_n534_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n598_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n600_), .A2(new_n602_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n590_), .B(new_n592_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n589_), .A3(new_n588_), .A4(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT37), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n609_), .A3(KEYINPUT37), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n503_), .B(new_n549_), .Z(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT16), .ZN(new_n621_));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(KEYINPUT17), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n618_), .B2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT72), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n614_), .A2(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n517_), .A2(new_n584_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n498_), .A3(new_n367_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n610_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n491_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n516_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n584_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n628_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n367_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G1gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n631_), .A2(new_n632_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n633_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n451_), .A2(new_n452_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n630_), .A2(new_n499_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n635_), .A2(new_n647_), .A3(new_n638_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G8gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G8gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT102), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(new_n648_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  AOI21_X1  g459(.A(new_n261_), .B1(new_n639_), .B2(new_n265_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n630_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n639_), .B2(new_n338_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT42), .Z(new_n667_));
  NAND3_X1  g466(.A1(new_n630_), .A2(new_n665_), .A3(new_n338_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n627_), .A2(new_n610_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT104), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n517_), .A2(new_n584_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n367_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n674_));
  INV_X1    g473(.A(new_n613_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT37), .B1(new_n606_), .B2(new_n609_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n491_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n457_), .A2(new_n463_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n487_), .B1(new_n484_), .B2(new_n339_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n265_), .B1(new_n682_), .B2(new_n488_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n679_), .B(new_n614_), .C1(new_n683_), .C2(new_n453_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n678_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n637_), .A2(new_n627_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n674_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(KEYINPUT44), .B2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n367_), .A2(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n673_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n672_), .A2(new_n692_), .A3(new_n647_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT45), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n689_), .A2(new_n647_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n694_), .B(new_n695_), .C1(new_n696_), .C2(new_n692_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n695_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n692_), .B1(new_n689_), .B2(new_n647_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n693_), .B(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n697_), .A2(new_n702_), .ZN(G1329gat));
  NAND3_X1  g502(.A1(new_n689_), .A2(G43gat), .A3(new_n265_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n672_), .A2(new_n265_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n256_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n709_), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n672_), .B2(new_n338_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n338_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n689_), .B2(new_n713_), .ZN(G1331gat));
  NOR3_X1   g513(.A1(new_n491_), .A2(new_n636_), .A3(new_n584_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n629_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n367_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n584_), .A2(new_n636_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n635_), .A2(new_n627_), .A3(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(new_n367_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n721_), .B2(new_n717_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n716_), .A2(new_n723_), .A3(new_n647_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n720_), .A2(new_n647_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G64gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT48), .B(new_n723_), .C1(new_n720_), .C2(new_n647_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n720_), .B2(new_n265_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT49), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n716_), .A2(new_n731_), .A3(new_n265_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1334gat));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n720_), .B2(new_n338_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n736_), .A3(new_n338_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  OR2_X1    g540(.A1(new_n685_), .A2(KEYINPUT108), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n685_), .A2(KEYINPUT108), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n719_), .A2(new_n628_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n368_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n715_), .A2(new_n671_), .ZN(new_n748_));
  INV_X1    g547(.A(G85gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n367_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1336gat));
  AOI21_X1  g550(.A(G92gat), .B1(new_n748_), .B2(new_n647_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n746_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n647_), .A2(new_n531_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT109), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n752_), .B1(new_n753_), .B2(new_n755_), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n746_), .B2(new_n490_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n715_), .A2(new_n265_), .A3(new_n526_), .A4(new_n671_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT110), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n757_), .B(new_n759_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n719_), .A2(new_n338_), .A3(new_n628_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n488_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n769_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n770_), .A2(new_n265_), .B1(new_n647_), .B2(new_n369_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n679_), .B1(new_n771_), .B2(new_n614_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n491_), .A2(KEYINPUT43), .A3(new_n677_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n527_), .B1(new_n685_), .B2(new_n768_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n775_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n767_), .B1(new_n678_), .B2(new_n684_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n782_), .C2(new_n527_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(KEYINPUT112), .A3(new_n775_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n778_), .A2(new_n781_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n748_), .A2(new_n527_), .A3(new_n338_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n789_), .A3(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n565_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n569_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(KEYINPUT55), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT114), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n793_), .A2(new_n794_), .A3(new_n797_), .A4(KEYINPUT55), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n552_), .ZN(new_n801_));
  OAI211_X1 g600(.A(G230gat), .B(G233gat), .C1(new_n565_), .C2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n796_), .A2(new_n798_), .A3(new_n800_), .A4(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n575_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT56), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(new_n806_), .A3(new_n575_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n507_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n504_), .A2(new_n506_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n515_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n809_), .B(new_n810_), .C1(new_n510_), .C2(new_n808_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n511_), .B2(new_n810_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n805_), .A2(new_n807_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n805_), .A2(KEYINPUT58), .A3(new_n807_), .A4(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n614_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n579_), .A2(new_n580_), .A3(new_n812_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n577_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n516_), .B1(new_n804_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n803_), .A2(new_n575_), .A3(new_n821_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n820_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n819_), .B1(new_n825_), .B2(new_n634_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n818_), .A2(new_n826_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n819_), .A3(new_n634_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n628_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n677_), .A2(new_n516_), .A3(new_n584_), .A4(new_n627_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT54), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n629_), .A2(new_n832_), .A3(new_n516_), .A4(new_n584_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n647_), .A2(new_n490_), .A3(new_n368_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n339_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n792_), .B1(new_n837_), .B2(new_n516_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n838_), .A2(KEYINPUT116), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(KEYINPUT116), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n338_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT59), .A3(new_n836_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n516_), .A2(new_n792_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n839_), .A2(new_n840_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(new_n837_), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n584_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n848_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n584_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n849_), .ZN(G1341gat));
  NAND2_X1  g652(.A1(new_n627_), .A2(KEYINPUT117), .ZN(new_n854_));
  MUX2_X1   g653(.A(KEYINPUT117), .B(new_n854_), .S(G127gat), .Z(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n844_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT59), .B1(new_n843_), .B2(new_n836_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n205_), .B1(new_n837_), .B2(new_n628_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n855_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n861_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1342gat));
  AOI21_X1  g665(.A(G134gat), .B1(new_n848_), .B2(new_n634_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT119), .B(G134gat), .Z(new_n868_));
  NOR2_X1   g667(.A1(new_n677_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n845_), .B2(new_n869_), .ZN(G1343gat));
  AOI21_X1  g669(.A(new_n265_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(new_n338_), .A3(new_n367_), .A4(new_n646_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n516_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n283_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n584_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n284_), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n872_), .A2(new_n628_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n872_), .B2(new_n677_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n634_), .A2(new_n273_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n872_), .B2(new_n881_), .ZN(G1347gat));
  INV_X1    g681(.A(new_n843_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n646_), .A2(new_n490_), .A3(new_n367_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n636_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT120), .ZN(new_n886_));
  OAI21_X1  g685(.A(G169gat), .B1(new_n883_), .B2(new_n886_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n843_), .A2(new_n890_), .A3(new_n884_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n843_), .B2(new_n884_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n636_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n888_), .A2(new_n889_), .B1(new_n894_), .B2(new_n895_), .ZN(G1348gat));
  NOR2_X1   g695(.A1(new_n584_), .A2(G176gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n835_), .A2(new_n339_), .A3(new_n884_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G176gat), .B1(new_n899_), .B2(new_n584_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n898_), .A2(KEYINPUT122), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902_));
  INV_X1    g701(.A(new_n897_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n899_), .A2(KEYINPUT121), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n891_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n900_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n902_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n901_), .A2(new_n907_), .ZN(G1349gat));
  NOR2_X1   g707(.A1(new_n628_), .A2(new_n416_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n237_), .B1(new_n899_), .B2(new_n628_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(KEYINPUT123), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  INV_X1    g712(.A(new_n909_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n904_), .B2(new_n891_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n911_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n913_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n912_), .A2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g717(.A(new_n634_), .B1(new_n243_), .B2(new_n381_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n677_), .B1(new_n904_), .B2(new_n891_), .ZN(new_n920_));
  INV_X1    g719(.A(G190gat), .ZN(new_n921_));
  OAI22_X1  g720(.A1(new_n894_), .A2(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n647_), .A2(new_n454_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n871_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n636_), .ZN(new_n927_));
  INV_X1    g726(.A(G197gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n926_), .A2(new_n931_), .A3(G197gat), .A4(new_n636_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n929_), .A2(new_n930_), .A3(new_n932_), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n925_), .A2(new_n584_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT125), .B(G204gat), .Z(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n934_), .B2(new_n937_), .ZN(G1353gat));
  NOR3_X1   g737(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n926_), .A2(new_n627_), .A3(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n941_), .B(new_n943_), .ZN(G1354gat));
  AND3_X1   g743(.A1(new_n926_), .A2(G218gat), .A3(new_n614_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n925_), .A2(new_n610_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n946_), .A2(KEYINPUT127), .ZN(new_n947_));
  AOI21_X1  g746(.A(G218gat), .B1(new_n946_), .B2(KEYINPUT127), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(G1355gat));
endmodule


