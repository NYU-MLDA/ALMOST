//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_;
  NAND2_X1  g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G57gat), .A2(G64gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT11), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G57gat), .ZN(new_n206_));
  INV_X1    g005(.A(G64gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(new_n202_), .ZN(new_n210_));
  INV_X1    g009(.A(G78gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G71gat), .ZN(new_n212_));
  INV_X1    g011(.A(G71gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G78gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n205_), .A2(new_n210_), .A3(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n209_), .B1(new_n208_), .B2(new_n202_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G85gat), .A3(G92gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT10), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(KEYINPUT10), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G85gat), .ZN(new_n233_));
  INV_X1    g032(.A(G92gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT9), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n229_), .A3(new_n228_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n240_), .A2(new_n222_), .A3(new_n225_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT8), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n235_), .A2(new_n236_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n219_), .B(new_n238_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G230gat), .ZN(new_n248_));
  INV_X1    g047(.A(G233gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n247_), .A2(KEYINPUT67), .A3(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n216_), .A2(new_n218_), .A3(KEYINPUT12), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT10), .B(G99gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n237_), .B1(new_n258_), .B2(G106gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT65), .B1(new_n259_), .B2(new_n226_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n227_), .A2(new_n232_), .A3(new_n261_), .A4(new_n237_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n242_), .A2(new_n244_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT8), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n263_), .A2(KEYINPUT66), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(new_n263_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n257_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n219_), .B1(new_n267_), .B2(new_n238_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT12), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n256_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n247_), .B(KEYINPUT64), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n250_), .B1(new_n274_), .B2(new_n271_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT69), .B(G120gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n273_), .A2(new_n275_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n273_), .A2(new_n275_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n281_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n289_), .B2(new_n282_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT13), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G71gat), .B(G99gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT79), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n296_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G190gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT76), .B(G190gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n302_), .B(new_n303_), .C1(new_n304_), .C2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT23), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(KEYINPUT77), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(G169gat), .B2(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT24), .A4(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n305_), .A2(new_n307_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n308_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT22), .B1(new_n308_), .B2(KEYINPUT78), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n309_), .A3(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n304_), .A2(G183gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n306_), .B(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n321_), .B(new_n316_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT30), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n300_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n328_), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(G120gat), .ZN(new_n332_));
  INV_X1    g131(.A(G127gat), .ZN(new_n333_));
  INV_X1    g132(.A(G134gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G113gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G127gat), .A2(G134gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n332_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(G120gat), .A3(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT31), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n331_), .B(new_n347_), .Z(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  OR2_X1    g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n353_), .A2(new_n354_), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n355_));
  NAND3_X1  g154(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  OAI22_X1  g161(.A1(KEYINPUT83), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n351_), .B(new_n352_), .C1(new_n357_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n351_), .B2(KEYINPUT1), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n351_), .A2(KEYINPUT1), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT1), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(KEYINPUT82), .A3(G155gat), .A4(G162gat), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n352_), .A4(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n361_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n353_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n344_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n365_), .A2(new_n343_), .A3(new_n341_), .A4(new_n373_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(KEYINPUT94), .A3(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n365_), .A2(new_n373_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n343_), .A4(new_n341_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n350_), .B(new_n377_), .C1(new_n383_), .C2(new_n376_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n349_), .A3(new_n382_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n386_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n348_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G197gat), .A2(G204gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT85), .B(G204gat), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT21), .B(new_n396_), .C1(new_n397_), .C2(G197gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399_));
  INV_X1    g198(.A(G197gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G204gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n398_), .B(new_n399_), .C1(new_n402_), .C2(KEYINPUT21), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n404_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n402_), .A3(KEYINPUT21), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n380_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT87), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n412_), .B(new_n408_), .C1(new_n380_), .C2(new_n409_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT84), .B(G233gat), .Z(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n411_), .A2(G228gat), .A3(new_n413_), .A4(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(G228gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(KEYINPUT87), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT88), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n423_), .A3(new_n418_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT89), .B1(new_n419_), .B2(new_n421_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n380_), .A2(new_n409_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G22gat), .B(G50gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT28), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n427_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n425_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n422_), .A2(KEYINPUT89), .A3(new_n424_), .A4(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G8gat), .B(G36gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT99), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(KEYINPUT99), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT90), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT19), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT22), .B(G169gat), .Z(new_n447_));
  NOR2_X1   g246(.A1(G183gat), .A2(G190gat), .ZN(new_n448_));
  OAI221_X1 g247(.A(new_n316_), .B1(new_n447_), .B2(G176gat), .C1(new_n324_), .C2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT26), .B(G190gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n303_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n315_), .A2(new_n451_), .A3(new_n307_), .A4(new_n317_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n453_), .A2(KEYINPUT98), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(KEYINPUT98), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n403_), .A3(new_n407_), .A4(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n408_), .B2(new_n326_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n446_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n408_), .A2(new_n453_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n403_), .A2(new_n318_), .A3(new_n407_), .A4(new_n325_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(KEYINPUT20), .A3(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n446_), .B(KEYINPUT91), .Z(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n442_), .B(new_n443_), .C1(new_n459_), .C2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n458_), .B(new_n446_), .C1(new_n408_), .C2(new_n453_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT92), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT92), .B1(new_n462_), .B2(new_n463_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n441_), .B(new_n466_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n465_), .A2(KEYINPUT27), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n440_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT27), .B1(new_n472_), .B2(new_n469_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n435_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n395_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n391_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n377_), .B1(new_n383_), .B2(new_n376_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n349_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n383_), .A2(KEYINPUT96), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n379_), .A2(new_n483_), .A3(new_n382_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n350_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n391_), .A3(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n472_), .A2(new_n469_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT97), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n479_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n490_));
  AOI211_X1 g289(.A(KEYINPUT33), .B(new_n391_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n472_), .A2(new_n486_), .A3(new_n469_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT97), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n441_), .A2(KEYINPUT32), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n466_), .B(new_n495_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n459_), .A2(new_n464_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n393_), .B(new_n496_), .C1(new_n497_), .C2(new_n495_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n489_), .A2(new_n494_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n435_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n393_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n474_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n474_), .A3(new_n501_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n348_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n476_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G29gat), .B(G36gat), .ZN(new_n509_));
  INV_X1    g308(.A(G43gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G50gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n509_), .B(G43gat), .ZN(new_n513_));
  INV_X1    g312(.A(G50gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n512_), .A2(new_n515_), .A3(KEYINPUT15), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT72), .B(G22gat), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(G15gat), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  INV_X1    g322(.A(G8gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT72), .B(G22gat), .ZN(new_n526_));
  INV_X1    g325(.A(G15gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n522_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G8gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n532_), .B(new_n533_), .C1(new_n516_), .C2(new_n531_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n531_), .B(new_n516_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G229gat), .A3(G233gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n308_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n400_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n534_), .A2(new_n536_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT101), .B1(new_n508_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT101), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n502_), .A2(new_n501_), .A3(new_n474_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(new_n503_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n348_), .B1(new_n549_), .B2(new_n500_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n547_), .B(new_n544_), .C1(new_n550_), .C2(new_n476_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n293_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n531_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(new_n219_), .Z(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G155gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT74), .B(G127gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT17), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n555_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n555_), .A2(KEYINPUT17), .A3(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT75), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n567_), .B2(new_n563_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G134gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(G162gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  INV_X1    g374(.A(new_n269_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n263_), .A2(new_n267_), .A3(KEYINPUT66), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n576_), .A2(new_n577_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n267_), .A2(new_n238_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n516_), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT35), .B(new_n575_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n520_), .B1(new_n269_), .B2(new_n268_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n584_));
  INV_X1    g383(.A(new_n580_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n573_), .B1(new_n587_), .B2(KEYINPUT71), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT36), .A3(new_n572_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n590_));
  INV_X1    g389(.A(new_n573_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n581_), .A2(new_n586_), .A3(new_n590_), .A4(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT37), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n569_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n552_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n523_), .A3(new_n393_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n292_), .A2(new_n544_), .A3(new_n568_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT102), .ZN(new_n601_));
  INV_X1    g400(.A(new_n508_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n593_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n394_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n598_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  INV_X1    g406(.A(new_n474_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n596_), .A2(new_n524_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT103), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n596_), .A2(new_n611_), .A3(new_n524_), .A4(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n604_), .B2(new_n474_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(KEYINPUT40), .A3(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1325gat));
  OAI21_X1  g420(.A(G15gat), .B1(new_n604_), .B2(new_n507_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT41), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n596_), .A2(new_n527_), .A3(new_n348_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  OAI21_X1  g424(.A(G22gat), .B1(new_n604_), .B2(new_n435_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT105), .Z(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(KEYINPUT42), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(KEYINPUT42), .ZN(new_n629_));
  INV_X1    g428(.A(new_n596_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n435_), .A2(G22gat), .ZN(new_n631_));
  OAI22_X1  g430(.A1(new_n628_), .A2(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n633_));
  INV_X1    g432(.A(new_n594_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n508_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n636_), .B(new_n594_), .C1(new_n550_), .C2(new_n476_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n292_), .A2(new_n544_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n640_), .A3(new_n569_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n633_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n639_), .B(new_n568_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n642_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n393_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n646_), .A2(KEYINPUT107), .A3(new_n393_), .A4(new_n647_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(G29gat), .A3(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n568_), .A2(new_n603_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n293_), .B(new_n654_), .C1(new_n546_), .C2(new_n551_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n393_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n474_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n646_), .B2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n552_), .A2(new_n662_), .A3(new_n608_), .A4(new_n653_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT45), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n655_), .A2(new_n667_), .A3(new_n662_), .A4(new_n608_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n659_), .A2(new_n660_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n661_), .B1(new_n664_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n661_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n666_), .A2(new_n668_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n608_), .B1(new_n644_), .B2(KEYINPUT44), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n673_), .B(new_n674_), .C1(new_n676_), .C2(new_n662_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n672_), .A2(new_n677_), .ZN(G1329gat));
  NAND4_X1  g477(.A1(new_n646_), .A2(G43gat), .A3(new_n348_), .A4(new_n647_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT109), .B(G43gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n655_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n507_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n655_), .B2(new_n434_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n646_), .A2(new_n434_), .A3(new_n647_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g489(.A1(new_n508_), .A2(new_n544_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(new_n603_), .A3(new_n293_), .A4(new_n568_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n206_), .A3(new_n394_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n691_), .B(KEYINPUT111), .Z(new_n694_));
  NAND2_X1  g493(.A1(new_n595_), .A2(new_n293_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT110), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT112), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n393_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n693_), .B1(new_n699_), .B2(new_n206_), .ZN(G1332gat));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n207_), .A3(new_n608_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G64gat), .B1(new_n692_), .B2(new_n474_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1333gat));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n213_), .A3(new_n348_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G71gat), .B1(new_n692_), .B2(new_n507_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT49), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1334gat));
  NAND3_X1  g507(.A1(new_n698_), .A2(new_n211_), .A3(new_n434_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G78gat), .B1(new_n692_), .B2(new_n435_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT50), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1335gat));
  NAND3_X1  g511(.A1(new_n694_), .A2(new_n293_), .A3(new_n653_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n233_), .B1(new_n713_), .B2(new_n394_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n568_), .A2(new_n544_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n638_), .A2(new_n293_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(G85gat), .A3(new_n393_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1336gat));
  OAI21_X1  g517(.A(new_n234_), .B1(new_n713_), .B2(new_n474_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(G92gat), .A3(new_n608_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1337gat));
  NOR3_X1   g520(.A1(new_n713_), .A2(new_n507_), .A3(new_n258_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n229_), .B1(new_n716_), .B2(new_n348_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n722_), .A2(KEYINPUT51), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT51), .B1(new_n722_), .B2(new_n723_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1338gat));
  NAND4_X1  g525(.A1(new_n638_), .A2(new_n434_), .A3(new_n293_), .A4(new_n715_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n434_), .A2(new_n228_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n729_), .A2(new_n730_), .B1(new_n713_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g532(.A1(new_n544_), .A2(new_n282_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n273_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT64), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n247_), .B(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n270_), .A2(new_n738_), .A3(new_n272_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n250_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n256_), .A2(new_n270_), .A3(KEYINPUT55), .A4(new_n272_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n288_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT56), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT113), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n746_), .B(KEYINPUT56), .C1(new_n742_), .C2(new_n288_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n743_), .A2(new_n744_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n734_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n535_), .A2(new_n533_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n532_), .B1(new_n516_), .B2(new_n531_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n752_), .B(new_n540_), .C1(new_n753_), .C2(new_n533_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(new_n543_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n286_), .B2(new_n290_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT114), .B(new_n755_), .C1(new_n286_), .C2(new_n290_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT57), .B(new_n603_), .C1(new_n751_), .C2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT116), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n603_), .B1(new_n751_), .B2(new_n760_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n742_), .B2(new_n288_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n282_), .B(new_n755_), .C1(new_n749_), .C2(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n594_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n745_), .A2(new_n747_), .A3(new_n749_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n758_), .B(new_n759_), .C1(new_n771_), .C2(new_n734_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(KEYINPUT57), .A4(new_n603_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n762_), .A2(new_n765_), .A3(new_n770_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n569_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n595_), .A2(new_n545_), .A3(new_n292_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n595_), .A2(new_n779_), .A3(new_n545_), .A4(new_n292_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n776_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n475_), .A2(new_n507_), .A3(new_n394_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n775_), .A2(KEYINPUT117), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n764_), .A2(new_n763_), .B1(new_n769_), .B2(new_n594_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n762_), .A4(new_n774_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n569_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n786_), .B1(new_n791_), .B2(new_n781_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n785_), .B1(new_n792_), .B2(new_n783_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n793_), .A2(new_n336_), .A3(new_n545_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n792_), .B2(new_n544_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1340gat));
  OAI211_X1 g595(.A(new_n293_), .B(new_n785_), .C1(new_n792_), .C2(new_n783_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G120gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n332_), .B1(new_n292_), .B2(KEYINPUT60), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n792_), .B(new_n799_), .C1(KEYINPUT60), .C2(new_n332_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(KEYINPUT118), .A3(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1341gat));
  NOR3_X1   g604(.A1(new_n793_), .A2(new_n333_), .A3(new_n569_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G127gat), .B1(new_n792_), .B2(new_n568_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1342gat));
  NOR3_X1   g607(.A1(new_n793_), .A2(new_n334_), .A3(new_n634_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G134gat), .B1(new_n792_), .B2(new_n593_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1343gat));
  AOI21_X1  g610(.A(new_n608_), .B1(new_n791_), .B2(new_n781_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n348_), .A2(new_n435_), .A3(new_n394_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n545_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(new_n360_), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n292_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n361_), .ZN(G1345gat));
  NOR2_X1   g617(.A1(new_n814_), .A2(new_n569_), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT61), .B(G155gat), .Z(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  NOR2_X1   g620(.A1(new_n814_), .A2(new_n603_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(G162gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n814_), .A2(new_n634_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(G162gat), .B2(new_n824_), .ZN(G1347gat));
  NOR2_X1   g624(.A1(new_n395_), .A2(new_n474_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n782_), .A2(new_n435_), .A3(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n545_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT62), .B1(new_n828_), .B2(new_n308_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(G169gat), .C1(new_n827_), .C2(new_n545_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n834_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT120), .B(KEYINPUT62), .C1(new_n828_), .C2(new_n308_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n831_), .A2(new_n835_), .A3(new_n836_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n447_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n775_), .A2(new_n569_), .B1(new_n780_), .B2(new_n778_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n434_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n842_), .B2(new_n826_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n826_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n841_), .A2(KEYINPUT121), .A3(new_n434_), .A4(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n839_), .B(new_n544_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n838_), .A2(new_n846_), .ZN(G1348gat));
  NAND2_X1  g646(.A1(new_n791_), .A2(new_n781_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(G176gat), .A3(new_n826_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n849_), .A2(new_n434_), .A3(new_n292_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n842_), .A2(new_n840_), .A3(new_n826_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n292_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OR3_X1    g652(.A1(new_n853_), .A2(KEYINPUT122), .A3(G176gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT122), .B1(new_n853_), .B2(G176gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n850_), .B1(new_n854_), .B2(new_n855_), .ZN(G1349gat));
  INV_X1    g655(.A(new_n303_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n568_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n858_));
  INV_X1    g657(.A(G183gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n827_), .B2(new_n569_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT123), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n858_), .A2(new_n863_), .A3(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1350gat));
  OAI211_X1 g664(.A(new_n450_), .B(new_n593_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n634_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n867_));
  INV_X1    g666(.A(G190gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n866_), .B(KEYINPUT124), .C1(new_n867_), .C2(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1351gat));
  AND2_X1   g672(.A1(new_n848_), .A2(new_n502_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n348_), .A2(new_n474_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n400_), .A3(new_n544_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G197gat), .B1(new_n876_), .B2(new_n545_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1352gat));
  NAND4_X1  g679(.A1(new_n848_), .A2(new_n502_), .A3(new_n293_), .A4(new_n875_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G204gat), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(KEYINPUT125), .A3(G204gat), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n884_), .B(new_n885_), .C1(new_n397_), .C2(new_n881_), .ZN(G1353gat));
  NAND3_X1  g685(.A1(new_n874_), .A2(new_n568_), .A3(new_n875_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT126), .Z(new_n891_));
  NAND2_X1  g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n888_), .A2(new_n889_), .A3(new_n891_), .A4(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n889_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n891_), .A2(new_n889_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n892_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n894_), .B(new_n895_), .C1(new_n887_), .C2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n876_), .A2(new_n899_), .A3(new_n634_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n877_), .A2(new_n593_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n899_), .B2(new_n901_), .ZN(G1355gat));
endmodule


