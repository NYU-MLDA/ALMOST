//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n969_, new_n970_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n203_), .A3(KEYINPUT21), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT26), .B(G190gat), .Z(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT25), .B(G183gat), .Z(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(new_n224_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(new_n212_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT92), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n220_), .B1(new_n234_), .B2(G176gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(KEYINPUT92), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n211_), .B(new_n227_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n223_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT83), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT83), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n221_), .A2(KEYINPUT81), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n221_), .A2(KEYINPUT81), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246_));
  INV_X1    g045(.A(G183gat), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT25), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n225_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT25), .B1(new_n246_), .B2(new_n247_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n244_), .A2(new_n245_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n242_), .A2(new_n243_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT22), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT84), .B1(new_n254_), .B2(G169gat), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n218_), .B(new_n255_), .C1(new_n233_), .C2(KEYINPUT84), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n220_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n211_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n259_));
  NOR3_X1   g058(.A1(new_n240_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT19), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n202_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n258_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n259_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n239_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT98), .A3(new_n262_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n227_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n211_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n252_), .A2(new_n211_), .A3(new_n257_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n263_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT99), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT99), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n272_), .A2(new_n276_), .A3(new_n263_), .A4(new_n273_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n264_), .A2(new_n268_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT18), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT101), .B1(new_n278_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n277_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n260_), .A2(new_n202_), .A3(new_n263_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT98), .B1(new_n267_), .B2(new_n262_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT101), .ZN(new_n288_));
  INV_X1    g087(.A(new_n282_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n272_), .A2(new_n273_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n262_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n237_), .A2(new_n238_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n293_), .A2(KEYINPUT93), .A3(new_n211_), .A4(new_n227_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT93), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n239_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n262_), .A2(new_n269_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n265_), .A2(new_n294_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n298_), .A3(new_n282_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT27), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n283_), .A2(new_n290_), .A3(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n292_), .A2(new_n298_), .A3(new_n282_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n282_), .B1(new_n292_), .B2(new_n298_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT27), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  OR2_X1    g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n310_));
  OR2_X1    g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n310_), .B(new_n311_), .C1(KEYINPUT1), .C2(new_n309_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT87), .B1(new_n309_), .B2(KEYINPUT1), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n307_), .B(new_n308_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n307_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G113gat), .B(G120gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(KEYINPUT86), .A3(new_n328_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n330_), .B(KEYINPUT4), .C1(new_n334_), .C2(new_n322_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n314_), .A2(new_n321_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(new_n332_), .A3(new_n340_), .A4(new_n333_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT94), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n330_), .B1(new_n334_), .B2(new_n322_), .ZN(new_n343_));
  OAI22_X1  g142(.A1(new_n338_), .A2(new_n342_), .B1(new_n343_), .B2(new_n337_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  OAI221_X1 g149(.A(new_n348_), .B1(new_n343_), .B2(new_n337_), .C1(new_n338_), .C2(new_n342_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT100), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT100), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n344_), .A2(new_n353_), .A3(new_n349_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT85), .B(G15gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  INV_X1    g157(.A(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT30), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n252_), .A2(new_n257_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n357_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n357_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G227gat), .ZN(new_n370_));
  INV_X1    g169(.A(G233gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n334_), .A2(KEYINPUT31), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT31), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n332_), .A2(new_n373_), .A3(new_n333_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n370_), .B(new_n371_), .C1(new_n372_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n370_), .A2(new_n371_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n369_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n375_), .A2(new_n378_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G78gat), .B(G106gat), .Z(new_n383_));
  XOR2_X1   g182(.A(G22gat), .B(G50gat), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n339_), .A2(KEYINPUT29), .A3(new_n386_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n383_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n394_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n339_), .A2(KEYINPUT29), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n397_), .B(KEYINPUT89), .Z(new_n398_));
  AND2_X1   g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n211_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n401_));
  OAI21_X1  g200(.A(new_n271_), .B1(new_n322_), .B2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n398_), .A2(new_n400_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n383_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n390_), .A2(new_n392_), .A3(KEYINPUT91), .A4(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n395_), .A2(new_n396_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n395_), .A2(new_n405_), .B1(new_n396_), .B2(new_n403_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n382_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n369_), .B(new_n380_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n395_), .A2(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n396_), .A2(new_n403_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n413_), .A3(new_n406_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n356_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n351_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n348_), .A2(KEYINPUT33), .ZN(new_n418_));
  OAI221_X1 g217(.A(new_n418_), .B1(new_n343_), .B2(new_n337_), .C1(new_n338_), .C2(new_n342_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n335_), .A2(new_n336_), .ZN(new_n420_));
  OAI221_X1 g219(.A(new_n349_), .B1(new_n343_), .B2(new_n336_), .C1(new_n420_), .C2(new_n342_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n292_), .A2(new_n298_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n289_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n299_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT96), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n421_), .A2(new_n419_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n304_), .A2(new_n427_), .A3(new_n428_), .A4(new_n417_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n282_), .A2(KEYINPUT32), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n278_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n352_), .B(new_n354_), .C1(new_n423_), .C2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n426_), .B(new_n429_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n410_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n306_), .A2(new_n415_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G229gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G29gat), .B(G36gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G43gat), .B(G50gat), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G43gat), .B(G50gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G8gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(G1gat), .ZN(new_n447_));
  INV_X1    g246(.A(G1gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G8gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT75), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n448_), .A2(KEYINPUT72), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT72), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G1gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n446_), .A2(KEYINPUT73), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G8gat), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n457_), .A2(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT14), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n456_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n457_), .A2(new_n459_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT73), .B(G8gat), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT74), .B(KEYINPUT14), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G15gat), .B(G22gat), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n455_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  AOI211_X1 g271(.A(new_n470_), .B(new_n454_), .C1(new_n465_), .C2(new_n468_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n445_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n457_), .A2(new_n459_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n460_), .A2(new_n462_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT74), .B1(new_n477_), .B2(KEYINPUT14), .ZN(new_n478_));
  AOI211_X1 g277(.A(new_n456_), .B(new_n464_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n471_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n454_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n469_), .A2(new_n471_), .A3(new_n455_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n445_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n474_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n474_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n438_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n442_), .A2(KEYINPUT15), .A3(new_n444_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT15), .B1(new_n442_), .B2(new_n444_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n481_), .A2(new_n491_), .A3(new_n482_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT79), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n481_), .A2(new_n491_), .A3(KEYINPUT79), .A4(new_n482_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n474_), .A3(new_n437_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n488_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT10), .B(G99gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(G106gat), .ZN(new_n510_));
  OR2_X1    g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n511_), .A2(KEYINPUT64), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT6), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(KEYINPUT9), .A3(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n524_), .A2(KEYINPUT9), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n520_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n515_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n520_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n523_), .A2(KEYINPUT65), .A3(new_n524_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n529_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  AOI211_X1 g336(.A(KEYINPUT8), .B(new_n535_), .C1(new_n533_), .C2(new_n520_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n528_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G64gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(G57gat), .ZN(new_n542_));
  INV_X1    g341(.A(G57gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(G64gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT11), .ZN(new_n548_));
  INV_X1    g347(.A(G78gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G71gat), .ZN(new_n550_));
  INV_X1    g349(.A(G71gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(G78gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n555_), .A2(KEYINPUT11), .A3(new_n542_), .A4(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n540_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n528_), .B(new_n557_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n507_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT67), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n548_), .A2(new_n553_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT11), .B1(new_n542_), .B2(new_n544_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n556_), .B(new_n562_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT12), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n562_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n515_), .A2(KEYINPUT66), .A3(new_n527_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT66), .B1(new_n515_), .B2(new_n527_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT68), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n540_), .B2(new_n557_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n568_), .B(new_n576_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n559_), .A2(new_n579_), .A3(new_n506_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n559_), .B2(new_n506_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n561_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT70), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(new_n590_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT13), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n584_), .A2(new_n590_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n595_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n540_), .B2(new_n445_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n491_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(KEYINPUT35), .B2(new_n603_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n607_), .A2(KEYINPUT35), .A3(new_n603_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n612_), .B(KEYINPUT36), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n609_), .B2(new_n614_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n616_), .A2(KEYINPUT37), .A3(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n619_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT17), .ZN(new_n628_));
  OAI211_X1 g427(.A(G231gat), .B(G233gat), .C1(new_n472_), .C2(new_n473_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n481_), .A2(new_n482_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(new_n557_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n557_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n628_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(KEYINPUT67), .A3(new_n635_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n632_), .A2(new_n557_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n562_), .B1(new_n638_), .B2(new_n633_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n627_), .A2(KEYINPUT17), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT77), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n636_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n622_), .A2(new_n643_), .ZN(new_n644_));
  NOR4_X1   g443(.A1(new_n436_), .A2(new_n505_), .A3(new_n599_), .A4(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n356_), .A3(new_n466_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n616_), .A2(new_n619_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n436_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n643_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n599_), .A2(new_n505_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n355_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n646_), .A2(new_n647_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n654_), .A3(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(new_n306_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n657_), .A3(new_n467_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n650_), .A2(KEYINPUT102), .A3(new_n657_), .A4(new_n652_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(G8gat), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n653_), .B2(new_n306_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n658_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n658_), .B(new_n667_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n653_), .B2(new_n382_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT41), .Z(new_n673_));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n645_), .A2(new_n674_), .A3(new_n410_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n407_), .A2(new_n408_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n645_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n653_), .B2(new_n678_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT104), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n436_), .A2(new_n505_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n651_), .A2(new_n649_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT106), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT106), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n599_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n686_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n356_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n599_), .A2(new_n505_), .A3(new_n643_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n426_), .A2(new_n429_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n433_), .A2(new_n431_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n435_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n409_), .A2(new_n414_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n700_), .A2(new_n301_), .A3(new_n305_), .A4(new_n355_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n622_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n696_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT43), .B(new_n622_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n694_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n694_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n356_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n693_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NOR2_X1   g511(.A1(new_n306_), .A2(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n686_), .A2(new_n690_), .A3(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n715_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n686_), .A2(new_n690_), .A3(new_n717_), .A4(new_n713_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n708_), .A2(new_n657_), .A3(new_n709_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G36gat), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n721_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1329gat));
  NOR2_X1   g527(.A1(new_n382_), .A2(new_n359_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n708_), .A2(new_n709_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n708_), .A2(KEYINPUT109), .A3(new_n709_), .A4(new_n729_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n359_), .B1(new_n691_), .B2(new_n382_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n733_), .A4(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n692_), .B2(new_n679_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n679_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n710_), .B2(new_n741_), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n643_), .A2(new_n505_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n650_), .A2(new_n599_), .A3(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n745_), .A2(new_n543_), .A3(new_n355_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  INV_X1    g546(.A(new_n505_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n436_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n702_), .A2(KEYINPUT110), .A3(new_n505_), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n598_), .B(new_n644_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT111), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT111), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n356_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n746_), .B1(new_n754_), .B2(new_n543_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n745_), .B2(new_n306_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  INV_X1    g556(.A(new_n751_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n657_), .A2(new_n541_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT112), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n758_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n745_), .B2(new_n382_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n751_), .A2(new_n551_), .A3(new_n410_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n745_), .B2(new_n678_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT113), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(KEYINPUT113), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(KEYINPUT50), .A3(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n751_), .A2(new_n549_), .A3(new_n679_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT50), .B1(new_n767_), .B2(new_n768_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n749_), .A2(new_n750_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n598_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n521_), .A3(new_n356_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n598_), .A2(new_n748_), .A3(new_n643_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n695_), .B1(new_n436_), .B2(new_n622_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n702_), .A2(new_n781_), .A3(new_n703_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n355_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n777_), .A2(new_n785_), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n776_), .A2(new_n522_), .A3(new_n657_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G92gat), .B1(new_n784_), .B2(new_n306_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1337gat));
  NOR2_X1   g588(.A1(new_n382_), .A2(new_n509_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n776_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT114), .ZN(new_n792_));
  INV_X1    g591(.A(G99gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n783_), .B2(new_n410_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n792_), .A2(KEYINPUT51), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT51), .B1(new_n792_), .B2(new_n794_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1338gat));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n780_), .A2(new_n782_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .A3(new_n679_), .A4(new_n778_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G106gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT116), .B1(new_n783_), .B2(new_n679_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n679_), .A3(new_n778_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(new_n800_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n678_), .A2(G106gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n774_), .A2(new_n775_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT115), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n774_), .A2(new_n811_), .A3(new_n775_), .A4(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n803_), .A2(new_n807_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT53), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n803_), .A2(new_n807_), .A3(new_n816_), .A4(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n575_), .A2(new_n577_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n559_), .A2(new_n506_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT69), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n580_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n822_), .A2(KEYINPUT55), .A3(new_n573_), .A4(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n573_), .A2(new_n577_), .A3(new_n575_), .A4(new_n559_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n507_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n821_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n588_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n474_), .A2(new_n438_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n501_), .B1(new_n496_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n437_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n588_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n561_), .B(new_n839_), .C1(new_n578_), .C2(new_n583_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n504_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n504_), .A2(new_n838_), .A3(KEYINPUT119), .A4(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n834_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n834_), .B2(new_n845_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n703_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n595_), .A2(new_n591_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n504_), .A2(new_n838_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n588_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT118), .ZN(new_n857_));
  INV_X1    g656(.A(new_n840_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n832_), .A2(new_n861_), .A3(new_n833_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n855_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n852_), .B1(new_n863_), .B2(new_n649_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n862_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n857_), .A2(new_n859_), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n865_), .A2(new_n866_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n649_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(KEYINPUT57), .A3(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n703_), .B(KEYINPUT120), .C1(new_n847_), .C2(new_n848_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n851_), .A2(new_n864_), .A3(new_n869_), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n651_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n853_), .A2(KEYINPUT13), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n596_), .B1(new_n595_), .B2(new_n591_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n643_), .A3(new_n505_), .A4(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n622_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT117), .B1(new_n744_), .B2(new_n598_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n744_), .A2(KEYINPUT117), .A3(new_n598_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n876_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .A4(new_n622_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n872_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n657_), .A2(new_n355_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n414_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n819_), .B1(new_n890_), .B2(new_n505_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT121), .B(new_n819_), .C1(new_n890_), .C2(new_n505_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n864_), .A2(new_n869_), .A3(new_n849_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n651_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n884_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n888_), .A2(KEYINPUT59), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n890_), .A2(KEYINPUT59), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n505_), .A2(new_n819_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n893_), .A2(new_n894_), .B1(new_n899_), .B2(new_n900_), .ZN(G1340gat));
  NAND2_X1  g700(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n898_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n599_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G120gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n888_), .B1(new_n872_), .B2(new_n884_), .ZN(new_n906_));
  INV_X1    g705(.A(G120gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n906_), .B(new_n908_), .C1(KEYINPUT60), .C2(new_n907_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n909_), .ZN(G1341gat));
  NAND3_X1  g709(.A1(new_n902_), .A2(new_n643_), .A3(new_n903_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G127gat), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n890_), .A2(G127gat), .A3(new_n651_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1342gat));
  INV_X1    g713(.A(G134gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n622_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n903_), .B(new_n916_), .C1(new_n906_), .C2(new_n917_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n843_), .A2(new_n844_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n856_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT58), .B1(new_n919_), .B2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n834_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT120), .B1(new_n924_), .B2(new_n703_), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n850_), .B(new_n622_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n863_), .A2(new_n852_), .A3(new_n649_), .ZN(new_n928_));
  AOI21_X1  g727(.A(KEYINPUT57), .B1(new_n867_), .B2(new_n868_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n643_), .B1(new_n927_), .B2(new_n930_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n879_), .A2(new_n883_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n649_), .B(new_n889_), .C1(new_n931_), .C2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n915_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n918_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n918_), .A2(new_n934_), .A3(KEYINPUT122), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1343gat));
  AOI21_X1  g738(.A(new_n932_), .B1(new_n871_), .B2(new_n651_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n409_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n941_), .A2(new_n748_), .A3(new_n886_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n599_), .A3(new_n886_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g744(.A1(new_n941_), .A2(new_n643_), .A3(new_n886_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT61), .B(G155gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n946_), .B(new_n947_), .ZN(G1346gat));
  NAND2_X1  g747(.A1(new_n941_), .A2(new_n886_), .ZN(new_n949_));
  OAI21_X1  g748(.A(G162gat), .B1(new_n949_), .B2(new_n622_), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n868_), .A2(G162gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n949_), .B2(new_n951_), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n306_), .A2(new_n356_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n414_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n897_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n748_), .ZN(new_n958_));
  XOR2_X1   g757(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n958_), .A2(G169gat), .A3(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n956_), .A2(new_n505_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n959_), .B1(new_n962_), .B2(new_n217_), .ZN(new_n963_));
  OAI211_X1 g762(.A(new_n961_), .B(new_n963_), .C1(new_n234_), .C2(new_n958_), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n957_), .B2(new_n599_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n940_), .A2(new_n679_), .ZN(new_n966_));
  NOR4_X1   g765(.A1(new_n954_), .A2(new_n218_), .A3(new_n382_), .A4(new_n598_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1349gat));
  NAND4_X1  g767(.A1(new_n966_), .A2(new_n410_), .A3(new_n643_), .A4(new_n953_), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n643_), .A2(new_n226_), .ZN(new_n970_));
  AOI22_X1  g769(.A1(new_n969_), .A2(new_n247_), .B1(new_n957_), .B2(new_n970_), .ZN(G1350gat));
  OAI21_X1  g770(.A(G190gat), .B1(new_n956_), .B2(new_n622_), .ZN(new_n972_));
  OR2_X1    g771(.A1(new_n868_), .A2(new_n225_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n956_), .B2(new_n973_), .ZN(G1351gat));
  NOR3_X1   g773(.A1(new_n940_), .A2(new_n409_), .A3(new_n954_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n748_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n599_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g778(.A(new_n651_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n980_));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n981_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n982_));
  OR3_X1    g781(.A1(new_n981_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983_));
  AOI22_X1  g782(.A1(new_n975_), .A2(new_n980_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n984_));
  AND2_X1   g783(.A1(new_n975_), .A2(new_n980_), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n984_), .B1(new_n985_), .B2(new_n983_), .ZN(G1354gat));
  INV_X1    g785(.A(new_n409_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(KEYINPUT125), .B(G218gat), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n703_), .A2(new_n988_), .ZN(new_n989_));
  XOR2_X1   g788(.A(new_n989_), .B(KEYINPUT126), .Z(new_n990_));
  NAND4_X1  g789(.A1(new_n885_), .A2(new_n987_), .A3(new_n953_), .A4(new_n990_), .ZN(new_n991_));
  NOR4_X1   g790(.A1(new_n940_), .A2(new_n409_), .A3(new_n868_), .A4(new_n954_), .ZN(new_n992_));
  OAI21_X1  g791(.A(new_n991_), .B1(new_n992_), .B2(new_n988_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n993_), .A2(KEYINPUT127), .ZN(new_n994_));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995_));
  OAI211_X1 g794(.A(new_n995_), .B(new_n991_), .C1(new_n992_), .C2(new_n988_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n994_), .A2(new_n996_), .ZN(G1355gat));
endmodule


