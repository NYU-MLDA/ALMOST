//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G64gat), .B(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  MUX2_X1   g012(.A(new_n212_), .B(KEYINPUT24), .S(new_n213_), .Z(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT76), .B(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT77), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n219_), .A2(KEYINPUT76), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(KEYINPUT76), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(KEYINPUT25), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(KEYINPUT78), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G190gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT79), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n230_), .B2(G190gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n227_), .B(new_n229_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n209_), .B(new_n214_), .C1(new_n223_), .C2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n210_), .A2(new_n211_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G169gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(new_n211_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n208_), .A2(new_n240_), .A3(KEYINPUT23), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n209_), .B2(new_n240_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n215_), .A2(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n239_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n236_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G197gat), .B(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT21), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G204gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G197gat), .ZN(new_n250_));
  INV_X1    g049(.A(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G204gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n252_), .A3(new_n247_), .ZN(new_n253_));
  AND2_X1   g052(.A1(G211gat), .A2(G218gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G211gat), .A2(G218gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n248_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n251_), .A2(G204gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n249_), .A2(G197gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n250_), .A2(new_n252_), .A3(KEYINPUT21), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n256_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n260_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI211_X1 g067(.A(KEYINPUT90), .B(new_n256_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n259_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(KEYINPUT92), .B(new_n259_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n245_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT19), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n239_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n229_), .A2(new_n231_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n281_), .B(new_n241_), .C1(new_n209_), .C2(new_n240_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n214_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n278_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n284_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n274_), .A2(new_n276_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n276_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n272_), .A2(new_n245_), .A3(new_n273_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT20), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n270_), .B2(new_n284_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n287_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n207_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n276_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n207_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n236_), .A2(new_n244_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n250_), .A2(new_n252_), .A3(KEYINPUT21), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT21), .B1(new_n250_), .B2(new_n252_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n267_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT90), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n266_), .A2(new_n260_), .A3(new_n267_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n258_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(KEYINPUT92), .ZN(new_n304_));
  AOI211_X1 g103(.A(new_n271_), .B(new_n258_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n297_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n285_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n287_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n295_), .A2(new_n296_), .A3(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n292_), .A2(new_n293_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n294_), .A2(new_n287_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n276_), .A3(new_n307_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n207_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT99), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT99), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n311_), .A2(new_n315_), .A3(new_n207_), .A4(new_n312_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n310_), .B1(new_n317_), .B2(KEYINPUT27), .ZN(new_n318_));
  XOR2_X1   g117(.A(G78gat), .B(G106gat), .Z(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(KEYINPUT94), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  AND2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  XOR2_X1   g130(.A(G141gat), .B(G148gat), .Z(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n339_), .A2(new_n342_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n323_), .A2(new_n322_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n335_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n335_), .A3(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI22_X1  g148(.A1(new_n333_), .A2(new_n334_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n303_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n321_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n330_), .A2(new_n332_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT86), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n345_), .A2(new_n346_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT87), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n348_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n355_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(KEYINPUT93), .B(new_n354_), .C1(new_n363_), .C2(new_n303_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n350_), .A2(KEYINPUT29), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n352_), .B(KEYINPUT89), .Z(new_n366_));
  OAI211_X1 g165(.A(new_n365_), .B(new_n366_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n353_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n319_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n353_), .A2(new_n364_), .A3(new_n367_), .A4(new_n319_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n320_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n373_));
  OR3_X1    g172(.A1(new_n350_), .A2(KEYINPUT29), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT94), .B1(new_n377_), .B2(new_n378_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n202_), .B1(new_n318_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(new_n371_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n386_), .A2(new_n381_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n316_), .A2(new_n309_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n293_), .B1(new_n388_), .B2(new_n314_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n387_), .B(KEYINPUT100), .C1(new_n389_), .C2(new_n310_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G127gat), .A2(G134gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(G113gat), .A2(G120gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G127gat), .A2(G134gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G113gat), .A2(G120gat), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(G127gat), .A2(G134gat), .ZN(new_n397_));
  AND2_X1   g196(.A1(G113gat), .A2(G120gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G113gat), .A2(G120gat), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n391_), .A2(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n396_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n362_), .B(new_n404_), .C1(new_n334_), .C2(new_n333_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n357_), .A2(new_n358_), .B1(new_n361_), .B2(new_n348_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n400_), .A2(KEYINPUT82), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n400_), .B2(KEYINPUT82), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n396_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n400_), .A2(KEYINPUT82), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT83), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n400_), .A2(KEYINPUT82), .A3(new_n407_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n396_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n405_), .B1(new_n406_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT4), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n410_), .A2(new_n415_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n350_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n417_), .A2(new_n419_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT0), .B(G57gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G85gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  NOR2_X1   g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n426_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n431_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n297_), .B(KEYINPUT30), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n438_), .A2(G43gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(G43gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G15gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(G71gat), .B(G99gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n439_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT81), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n445_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n448_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n447_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n384_), .A2(new_n390_), .A3(new_n437_), .A4(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n296_), .A2(KEYINPUT32), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n295_), .A2(new_n308_), .A3(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n274_), .A2(new_n287_), .A3(new_n285_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n276_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT32), .A3(new_n296_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n458_), .B(new_n462_), .C1(new_n432_), .C2(new_n435_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n286_), .A2(new_n291_), .A3(new_n207_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n296_), .B1(new_n295_), .B2(new_n308_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT96), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT96), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n292_), .A2(new_n309_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n427_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n433_), .A2(KEYINPUT33), .A3(new_n434_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n466_), .A2(new_n468_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n422_), .A2(new_n420_), .A3(new_n405_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT4), .B1(new_n421_), .B2(new_n350_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(KEYINPUT4), .B2(new_n417_), .ZN(new_n475_));
  OAI211_X1 g274(.A(KEYINPUT98), .B(new_n473_), .C1(new_n475_), .C2(new_n420_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n418_), .A2(new_n424_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT98), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n419_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(KEYINPUT33), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n431_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n463_), .B1(new_n472_), .B2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n315_), .B1(new_n461_), .B2(new_n207_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n316_), .A2(new_n309_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT27), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n310_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n486_), .A2(new_n487_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n483_), .A2(new_n387_), .B1(new_n488_), .B2(new_n437_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n456_), .B1(new_n489_), .B2(new_n455_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G232gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT34), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G85gat), .B(G92gat), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT6), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT68), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT68), .B1(new_n499_), .B2(new_n501_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(KEYINPUT7), .ZN(new_n507_));
  NOR2_X1   g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n507_), .A2(new_n508_), .B1(new_n505_), .B2(KEYINPUT7), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT66), .B1(new_n510_), .B2(KEYINPUT67), .ZN(new_n511_));
  OR2_X1    g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n497_), .B1(new_n504_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n500_), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n498_), .A2(KEYINPUT6), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n509_), .A2(new_n519_), .A3(new_n513_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n496_), .A2(new_n516_), .ZN(new_n521_));
  OAI22_X1  g320(.A1(new_n515_), .A2(new_n516_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT9), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n496_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n519_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT10), .B(G99gat), .Z(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT64), .B(G106gat), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n524_), .A2(new_n525_), .A3(G85gat), .A4(G92gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n528_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G43gat), .ZN(new_n534_));
  OR2_X1    g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n539_));
  AOI21_X1  g338(.A(G50gat), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  INV_X1    g340(.A(G50gat), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n522_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n507_), .A2(new_n508_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n505_), .A2(KEYINPUT7), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT68), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n516_), .B1(new_n552_), .B2(new_n496_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n521_), .B1(new_n514_), .B2(new_n528_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n533_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT69), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT69), .B(new_n533_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT15), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n540_), .A2(new_n543_), .A3(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n542_), .B1(new_n541_), .B2(new_n537_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n538_), .A2(G50gat), .A3(new_n539_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT15), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT72), .B1(new_n559_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568_));
  AOI211_X1 g367(.A(new_n568_), .B(new_n565_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n495_), .B(new_n545_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n493_), .A2(new_n494_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT69), .B1(new_n522_), .B2(new_n533_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n558_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n566_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n568_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n559_), .A2(KEYINPUT72), .A3(new_n566_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n571_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n495_), .A4(new_n545_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n580_), .A3(KEYINPUT73), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G134gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G162gat), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n545_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n579_), .B1(new_n588_), .B2(new_n495_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n570_), .A2(new_n571_), .ZN(new_n590_));
  OAI211_X1 g389(.A(KEYINPUT36), .B(new_n584_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n585_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n572_), .A2(new_n580_), .A3(KEYINPUT73), .A4(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n586_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT37), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n586_), .A2(new_n591_), .A3(new_n596_), .A4(new_n593_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G15gat), .B(G22gat), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  INV_X1    g398(.A(G8gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT14), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G1gat), .B(G8gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  XNOR2_X1  g403(.A(G57gat), .B(G64gat), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT11), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(KEYINPUT11), .ZN(new_n607_));
  XOR2_X1   g406(.A(G71gat), .B(G78gat), .Z(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n604_), .B(new_n611_), .Z(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT16), .B(G183gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n614_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n620_), .B2(new_n614_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT74), .Z(new_n624_));
  AND3_X1   g423(.A1(new_n595_), .A2(new_n597_), .A3(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n555_), .A2(new_n610_), .A3(new_n609_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n533_), .B(new_n611_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(G230gat), .A3(G233gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT12), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n611_), .A2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n559_), .A2(new_n631_), .B1(new_n630_), .B2(new_n626_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT71), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT70), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n627_), .A2(KEYINPUT70), .A3(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n632_), .A2(new_n633_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n633_), .B1(new_n632_), .B2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n629_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(new_n249_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT5), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(new_n211_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n642_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n632_), .A2(new_n639_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT71), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n632_), .A2(new_n633_), .A3(new_n639_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n646_), .B1(new_n652_), .B2(new_n629_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT13), .B1(new_n648_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n642_), .A2(new_n647_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n629_), .A3(new_n646_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT13), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n654_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n544_), .A2(new_n604_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT75), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT75), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n544_), .A2(new_n604_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n544_), .B2(new_n604_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(G229gat), .A2(G233gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n565_), .A2(new_n604_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n666_), .A3(new_n664_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(new_n210_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(new_n251_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n668_), .A2(new_n670_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n659_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AND4_X1   g480(.A1(KEYINPUT101), .A2(new_n490_), .A3(new_n625_), .A4(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n455_), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n469_), .B(new_n431_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n292_), .A2(new_n309_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(KEYINPUT96), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(new_n481_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n383_), .B1(new_n687_), .B2(new_n463_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n318_), .A2(new_n387_), .A3(new_n436_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n683_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n680_), .B1(new_n690_), .B2(new_n456_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n691_), .B2(new_n625_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n682_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n436_), .B(KEYINPUT102), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n599_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n624_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n594_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n691_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G1gat), .B1(new_n700_), .B2(new_n437_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(KEYINPUT103), .A3(new_n696_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT103), .B1(new_n695_), .B2(new_n696_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n697_), .B(new_n701_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT104), .ZN(new_n706_));
  INV_X1    g505(.A(new_n704_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n702_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n697_), .A4(new_n701_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1324gat));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n693_), .A2(KEYINPUT105), .A3(new_n600_), .A4(new_n318_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n490_), .A2(new_n625_), .A3(new_n681_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n691_), .A2(KEYINPUT101), .A3(new_n625_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n600_), .A3(new_n318_), .A4(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n714_), .A2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n490_), .A2(new_n681_), .A3(new_n318_), .A4(new_n699_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT39), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G8gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G8gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n713_), .B1(new_n722_), .B2(new_n728_), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT106), .B(new_n727_), .C1(new_n714_), .C2(new_n721_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n712_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n719_), .A2(new_n720_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n719_), .A2(new_n720_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT106), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n722_), .A2(new_n713_), .A3(new_n728_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT40), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n731_), .A2(new_n737_), .ZN(G1325gat));
  OAI21_X1  g537(.A(G15gat), .B1(new_n700_), .B2(new_n683_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT41), .Z(new_n740_));
  INV_X1    g539(.A(new_n693_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n683_), .A2(G15gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(G1326gat));
  OAI21_X1  g542(.A(G22gat), .B1(new_n700_), .B2(new_n387_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT42), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n387_), .A2(G22gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n741_), .B2(new_n746_), .ZN(G1327gat));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n748_));
  INV_X1    g547(.A(new_n594_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n624_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n698_), .A2(KEYINPUT109), .A3(new_n594_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n691_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G29gat), .B1(new_n753_), .B2(new_n436_), .ZN(new_n754_));
  INV_X1    g553(.A(G29gat), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n680_), .A2(new_n624_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n595_), .A2(new_n597_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n490_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(KEYINPUT43), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n490_), .B2(new_n757_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT108), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(KEYINPUT108), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n758_), .A2(new_n760_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(KEYINPUT43), .B2(new_n758_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT108), .A3(new_n764_), .A4(new_n756_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n755_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n754_), .B1(new_n771_), .B2(new_n694_), .ZN(G1328gat));
  INV_X1    g571(.A(G36gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n753_), .A2(new_n773_), .A3(new_n318_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT45), .ZN(new_n775_));
  INV_X1    g574(.A(new_n318_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(new_n773_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1329gat));
  NAND3_X1  g579(.A1(new_n753_), .A2(new_n534_), .A3(new_n455_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n683_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n534_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(G1330gat));
  NAND2_X1  g584(.A1(new_n383_), .A2(new_n542_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT110), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n753_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n387_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n542_), .ZN(G1331gat));
  AOI211_X1 g589(.A(new_n679_), .B(new_n659_), .C1(new_n690_), .C2(new_n456_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n625_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT111), .Z(new_n793_));
  AOI21_X1  g592(.A(G57gat), .B1(new_n793_), .B2(new_n694_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n791_), .A2(G57gat), .A3(new_n436_), .A4(new_n699_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT112), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1332gat));
  NAND2_X1  g596(.A1(new_n791_), .A2(new_n699_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G64gat), .B1(new_n798_), .B2(new_n776_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT48), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n776_), .A2(G64gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT113), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n792_), .B2(new_n802_), .ZN(G1333gat));
  OAI21_X1  g602(.A(G71gat), .B1(new_n798_), .B2(new_n683_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT49), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n683_), .A2(G71gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n792_), .B2(new_n806_), .ZN(G1334gat));
  OAI21_X1  g606(.A(G78gat), .B1(new_n798_), .B2(new_n387_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT50), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n387_), .A2(G78gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n792_), .B2(new_n810_), .ZN(G1335gat));
  NOR3_X1   g610(.A1(new_n659_), .A2(new_n624_), .A3(new_n679_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n769_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G85gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n437_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n791_), .A2(new_n752_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G85gat), .B1(new_n817_), .B2(new_n694_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n815_), .A2(new_n818_), .ZN(G1336gat));
  NAND3_X1  g618(.A1(new_n769_), .A2(G92gat), .A3(new_n812_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n816_), .A2(new_n776_), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n820_), .A2(new_n776_), .B1(G92gat), .B2(new_n821_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT114), .Z(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n813_), .B2(new_n683_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n529_), .A3(new_n455_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n826_), .B(new_n827_), .Z(G1338gat));
  OAI211_X1 g627(.A(new_n383_), .B(new_n812_), .C1(new_n759_), .C2(new_n762_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G106gat), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT116), .A3(G106gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(KEYINPUT52), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n817_), .A2(new_n530_), .A3(new_n383_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n831_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT53), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n834_), .A2(new_n840_), .A3(new_n835_), .A4(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1339gat));
  XNOR2_X1  g641(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n625_), .A2(new_n678_), .A3(new_n659_), .A4(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n595_), .A2(new_n659_), .A3(new_n597_), .A4(new_n624_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n846_), .B2(new_n679_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n648_), .A2(new_n678_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n632_), .A2(KEYINPUT55), .A3(new_n639_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n634_), .B1(new_n632_), .B2(new_n627_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT56), .B1(new_n855_), .B2(new_n647_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n857_), .B(new_n646_), .C1(new_n851_), .C2(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n849_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n665_), .A2(new_n666_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n669_), .A2(new_n667_), .A3(new_n664_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n673_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n675_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n675_), .B2(new_n862_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n594_), .B1(new_n859_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT57), .B1(new_n869_), .B2(KEYINPUT119), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(new_n650_), .B2(new_n651_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n632_), .A2(new_n627_), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n874_), .A2(new_n634_), .B1(new_n850_), .B2(new_n649_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n647_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n857_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n855_), .A2(KEYINPUT56), .A3(new_n647_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n867_), .B1(new_n879_), .B2(new_n849_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n871_), .B(new_n872_), .C1(new_n880_), .C2(new_n594_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n866_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n656_), .B(new_n882_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n879_), .A2(KEYINPUT58), .A3(new_n656_), .A4(new_n882_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n757_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n870_), .A2(new_n881_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n848_), .B1(new_n698_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n694_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n384_), .A2(new_n390_), .A3(new_n455_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G113gat), .B1(new_n894_), .B2(new_n679_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n889_), .B2(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n888_), .A2(new_n698_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n848_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(KEYINPUT59), .A3(new_n892_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n678_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n895_), .B1(new_n902_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n659_), .B2(KEYINPUT60), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n894_), .B(new_n905_), .C1(KEYINPUT60), .C2(new_n904_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n659_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n904_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT120), .B(new_n906_), .C1(new_n907_), .C2(new_n904_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1341gat));
  AOI21_X1  g711(.A(G127gat), .B1(new_n894_), .B2(new_n624_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n698_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g714(.A(G134gat), .B1(new_n894_), .B2(new_n594_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n757_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n918_), .B2(G134gat), .ZN(G1343gat));
  NAND3_X1  g718(.A1(new_n900_), .A2(new_n683_), .A3(new_n383_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n694_), .A2(new_n776_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n920_), .A2(new_n678_), .A3(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT121), .B(G141gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1344gat));
  NOR2_X1   g723(.A1(new_n920_), .A2(new_n921_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n659_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g727(.A1(new_n925_), .A2(new_n624_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G155gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  AOI21_X1  g730(.A(G162gat), .B1(new_n925_), .B2(new_n594_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n920_), .A2(new_n917_), .A3(new_n921_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935_));
  NOR4_X1   g734(.A1(new_n694_), .A2(new_n683_), .A3(new_n776_), .A4(new_n383_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n900_), .A2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n937_), .B2(new_n678_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n900_), .A2(KEYINPUT122), .A3(new_n679_), .A4(new_n936_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n938_), .A2(G169gat), .A3(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n937_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n943_), .A2(new_n679_), .A3(new_n238_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n938_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n939_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n944_), .A3(new_n945_), .ZN(G1348gat));
  NOR2_X1   g745(.A1(new_n937_), .A2(new_n659_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n211_), .ZN(G1349gat));
  NOR2_X1   g747(.A1(new_n937_), .A2(new_n698_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n949_), .A2(new_n280_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n215_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n949_), .A2(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(KEYINPUT123), .B1(new_n950_), .B2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n949_), .A2(new_n280_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955_));
  OAI211_X1 g754(.A(new_n954_), .B(new_n955_), .C1(new_n951_), .C2(new_n949_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n953_), .A2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n937_), .B2(new_n917_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n958_), .B(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n943_), .A2(new_n594_), .A3(new_n279_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1351gat));
  NOR2_X1   g761(.A1(new_n776_), .A2(new_n436_), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n900_), .A2(new_n683_), .A3(new_n383_), .A4(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n678_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(new_n251_), .ZN(G1352gat));
  NOR3_X1   g765(.A1(new_n889_), .A2(new_n455_), .A3(new_n387_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n967_), .A2(new_n926_), .A3(new_n963_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(G204gat), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n970_), .B1(KEYINPUT125), .B2(new_n249_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n968_), .A2(new_n969_), .A3(G204gat), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(G1353gat));
  NOR2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n974_), .B1(new_n964_), .B2(new_n698_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(KEYINPUT126), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  OAI211_X1 g776(.A(new_n977_), .B(new_n974_), .C1(new_n964_), .C2(new_n698_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n964_), .A2(new_n698_), .ZN(new_n979_));
  XOR2_X1   g778(.A(KEYINPUT63), .B(G211gat), .Z(new_n980_));
  AOI22_X1  g779(.A1(new_n976_), .A2(new_n978_), .B1(new_n979_), .B2(new_n980_), .ZN(G1354gat));
  OAI21_X1  g780(.A(G218gat), .B1(new_n964_), .B2(new_n917_), .ZN(new_n982_));
  INV_X1    g781(.A(G218gat), .ZN(new_n983_));
  NAND4_X1  g782(.A1(new_n967_), .A2(new_n983_), .A3(new_n594_), .A4(new_n963_), .ZN(new_n984_));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n982_), .A2(new_n984_), .A3(new_n985_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n985_), .B1(new_n982_), .B2(new_n984_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1355gat));
endmodule


