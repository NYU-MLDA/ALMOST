//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT78), .B(KEYINPUT25), .ZN(new_n207_));
  OAI211_X1 g006(.A(KEYINPUT79), .B(new_n206_), .C1(new_n207_), .C2(new_n205_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n204_), .A2(KEYINPUT78), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n215_), .A3(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n208_), .A2(new_n212_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n221_), .A2(KEYINPUT81), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT81), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(KEYINPUT24), .A3(new_n230_), .ZN(new_n231_));
  OR3_X1    g030(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n219_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n221_), .A2(new_n224_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT22), .ZN(new_n237_));
  AOI21_X1  g036(.A(G176gat), .B1(new_n237_), .B2(KEYINPUT82), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G169gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n228_), .ZN(new_n240_));
  OAI221_X1 g039(.A(new_n236_), .B1(new_n227_), .B2(new_n238_), .C1(KEYINPUT82), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G211gat), .B(G218gat), .Z(new_n243_));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(G197gat), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n246_), .A2(new_n248_), .B1(G197gat), .B2(new_n245_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G197gat), .B(G204gat), .Z(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(KEYINPUT21), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n250_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n243_), .A2(new_n251_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n242_), .A2(new_n256_), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n222_), .A2(new_n225_), .B1(G183gat), .B2(G190gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n240_), .A2(new_n230_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n231_), .A2(new_n235_), .A3(new_n232_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT25), .B(G183gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n258_), .A2(new_n259_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT20), .B1(new_n264_), .B2(new_n255_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n203_), .B1(new_n257_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n242_), .A2(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n203_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n255_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n267_), .A2(KEYINPUT20), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT18), .B(G64gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G92gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n266_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G113gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT83), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G113gat), .ZN(new_n281_));
  INV_X1    g080(.A(G120gat), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G134gat), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n280_), .A2(G113gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n278_), .A2(KEYINPUT83), .ZN(new_n289_));
  OAI21_X1  g088(.A(G120gat), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n301_));
  NOR2_X1   g100(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n296_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT85), .B(new_n296_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n294_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n294_), .A2(KEYINPUT1), .ZN(new_n315_));
  INV_X1    g114(.A(new_n308_), .ZN(new_n316_));
  AND2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n317_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n293_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n286_), .A2(new_n292_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n312_), .B(new_n300_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(new_n294_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(KEYINPUT4), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT4), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n293_), .B(new_n326_), .C1(new_n314_), .C2(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT93), .Z(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n320_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n330_), .A2(KEYINPUT33), .A3(new_n331_), .A4(new_n335_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n277_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n325_), .A2(new_n328_), .A3(new_n327_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n335_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n320_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT94), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n341_), .A2(new_n346_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n340_), .A2(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n257_), .A2(new_n265_), .A3(new_n203_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n267_), .A2(KEYINPUT20), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n269_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n203_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n336_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n330_), .A2(KEYINPUT95), .A3(new_n331_), .A4(new_n335_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n330_), .A2(new_n331_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT96), .B1(new_n360_), .B2(new_n342_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT96), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n362_), .B(new_n335_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n355_), .B1(new_n359_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n266_), .A2(new_n270_), .A3(new_n354_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n349_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n307_), .A2(new_n313_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n294_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n319_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n256_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G228gat), .ZN(new_n375_));
  INV_X1    g174(.A(G233gat), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n376_), .A2(KEYINPUT88), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(KEYINPUT88), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT89), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n256_), .B(new_n380_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n372_), .A2(new_n373_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G22gat), .B(G50gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n388_));
  INV_X1    g187(.A(new_n386_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n372_), .A2(new_n373_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n388_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n389_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n393_));
  NOR4_X1   g192(.A1(new_n314_), .A2(new_n319_), .A3(KEYINPUT29), .A4(new_n386_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n369_), .B(new_n384_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n384_), .A2(new_n369_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n397_), .A3(new_n395_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT91), .B1(new_n391_), .B2(new_n395_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n382_), .A2(new_n368_), .A3(new_n383_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n399_), .B(new_n400_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n401_), .A2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n398_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT97), .B1(new_n367_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n360_), .A2(new_n342_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n362_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n360_), .A2(KEYINPUT96), .A3(new_n342_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n277_), .A2(KEYINPUT27), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n277_), .A2(KEYINPUT99), .A3(KEYINPUT27), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n275_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n274_), .B(KEYINPUT98), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n418_), .B(KEYINPUT27), .C1(new_n353_), .C2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n412_), .A2(new_n417_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n355_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n411_), .A2(new_n366_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n348_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(new_n277_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT97), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n407_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n406_), .A2(new_n421_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(new_n321_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G15gat), .B(G43gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT31), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n435_), .A2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n433_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n432_), .A3(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n429_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n411_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n420_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n448_), .A2(new_n405_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(G57gat), .A2(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G57gat), .A2(G64gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT11), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G78gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n459_), .A3(new_n454_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(new_n457_), .A3(KEYINPUT11), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G231gat), .A2(G233gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  AND2_X1   g264(.A1(G1gat), .A2(G8gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT14), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(G15gat), .A2(G22gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G15gat), .A2(G22gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OR3_X1    g270(.A1(new_n468_), .A2(new_n471_), .A3(KEYINPUT74), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G1gat), .A2(G8gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n466_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT74), .B1(new_n468_), .B2(new_n471_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n465_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G127gat), .B(G155gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G183gat), .B(G211gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n480_), .A2(new_n481_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(KEYINPUT17), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n480_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n452_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT10), .B(G99gat), .Z(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G85gat), .B(G92gat), .Z(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT9), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n497_));
  NOR2_X1   g296(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(G92gat), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n493_), .A2(new_n495_), .A3(new_n499_), .A4(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n492_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n508_), .A2(new_n502_), .A3(new_n503_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n494_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(KEYINPUT8), .A3(new_n494_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n463_), .A2(new_n505_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT66), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT12), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G230gat), .A2(G233gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n505_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n463_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n516_), .A2(KEYINPUT12), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n518_), .B(new_n519_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(KEYINPUT65), .A3(new_n515_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n528_), .A3(new_n521_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n525_), .B1(new_n530_), .B2(new_n519_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n245_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G176gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n531_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT67), .B(KEYINPUT13), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n539_), .B2(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G29gat), .B(G36gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n544_), .A2(new_n545_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n479_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n478_), .B1(new_n551_), .B2(new_n549_), .ZN(new_n554_));
  OAI211_X1 g353(.A(G229gat), .B(G233gat), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n551_), .A3(KEYINPUT15), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n550_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n542_), .B1(new_n550_), .B2(new_n546_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n478_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT76), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n479_), .A2(new_n552_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT77), .Z(new_n565_));
  INV_X1    g364(.A(KEYINPUT76), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n478_), .A2(new_n566_), .A3(new_n556_), .A4(new_n560_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .A4(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n227_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n247_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n555_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n555_), .B2(new_n568_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n541_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n490_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n560_), .A2(new_n556_), .A3(new_n520_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n552_), .A2(new_n505_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT68), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n580_), .B2(KEYINPUT71), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n582_), .A2(new_n586_), .B1(new_n588_), .B2(new_n585_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n582_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT72), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G134gat), .ZN(new_n593_));
  INV_X1    g392(.A(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT36), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n582_), .A2(new_n586_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n588_), .A2(new_n585_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n582_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n596_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n606_), .B(new_n595_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n591_), .A2(new_n602_), .A3(KEYINPUT73), .A4(new_n596_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n601_), .A3(new_n596_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n579_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(G1gat), .A3(new_n447_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n579_), .A2(new_n609_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n447_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(new_n489_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n578_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n449_), .A4(new_n609_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(new_n627_), .A3(G8gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n626_), .B2(G8gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n449_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(G8gat), .ZN(new_n631_));
  OAI22_X1  g430(.A1(new_n628_), .A2(new_n629_), .B1(new_n616_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT101), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634_));
  OAI221_X1 g433(.A(new_n634_), .B1(new_n616_), .B2(new_n631_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n633_), .A2(KEYINPUT40), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT40), .B1(new_n633_), .B2(new_n635_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1325gat));
  NOR3_X1   g437(.A1(new_n616_), .A2(G15gat), .A3(new_n445_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT102), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n579_), .A2(new_n444_), .A3(new_n609_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n641_), .B2(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  OAI21_X1  g443(.A(G22gat), .B1(new_n620_), .B2(new_n407_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n407_), .A2(G22gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n616_), .B2(new_n647_), .ZN(G1327gat));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n614_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n614_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n611_), .A2(KEYINPUT103), .A3(new_n613_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n427_), .B1(new_n426_), .B2(new_n407_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT97), .B(new_n405_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n444_), .B1(new_n659_), .B2(new_n421_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n660_), .B2(new_n450_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n652_), .B1(new_n661_), .B2(KEYINPUT43), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n578_), .A2(new_n489_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n649_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n650_), .B1(new_n452_), .B2(new_n656_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT44), .B(new_n663_), .C1(new_n666_), .C2(new_n652_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G29gat), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n447_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n450_), .B1(new_n429_), .B2(new_n445_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n609_), .A3(new_n664_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n411_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT104), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n665_), .A2(new_n449_), .A3(new_n667_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(KEYINPUT104), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n609_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n452_), .A2(new_n680_), .A3(new_n663_), .A4(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT45), .B1(new_n682_), .B2(new_n630_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n672_), .A2(new_n684_), .A3(new_n680_), .A4(new_n449_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  AND4_X1   g485(.A1(new_n676_), .A2(new_n678_), .A3(new_n679_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n686_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n677_), .B2(G36gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n676_), .B1(new_n689_), .B2(new_n679_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1329gat));
  NAND2_X1  g490(.A1(new_n444_), .A2(G43gat), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n672_), .A2(new_n444_), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n668_), .A2(new_n692_), .B1(G43gat), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n672_), .A2(new_n696_), .A3(new_n405_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n665_), .A2(new_n405_), .A3(new_n667_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n698_), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n698_), .B2(G50gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1331gat));
  INV_X1    g500(.A(G57gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n541_), .A2(new_n577_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n624_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n615_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n705_), .B2(new_n447_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n624_), .A2(new_n609_), .A3(new_n703_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n624_), .A2(KEYINPUT106), .A3(new_n609_), .A4(new_n703_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n709_), .A2(G57gat), .A3(new_n411_), .A4(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n706_), .A2(new_n711_), .ZN(G1332gat));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n449_), .A3(new_n710_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G64gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n630_), .A2(G64gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT107), .Z(new_n718_));
  OAI22_X1  g517(.A1(new_n715_), .A2(new_n716_), .B1(new_n705_), .B2(new_n718_), .ZN(G1333gat));
  OR3_X1    g518(.A1(new_n705_), .A2(G71gat), .A3(new_n445_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n709_), .A2(new_n444_), .A3(new_n710_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT49), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT108), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1334gat));
  OR3_X1    g528(.A1(new_n705_), .A2(G78gat), .A3(new_n407_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n709_), .A2(new_n405_), .A3(new_n710_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(G78gat), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G78gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT110), .B(new_n730_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1335gat));
  NOR3_X1   g538(.A1(new_n541_), .A2(new_n577_), .A3(new_n489_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n671_), .A2(new_n609_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n411_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n661_), .A2(KEYINPUT43), .ZN(new_n746_));
  INV_X1    g545(.A(new_n652_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT112), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n662_), .A2(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(new_n740_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n498_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n447_), .B1(new_n753_), .B2(new_n496_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n745_), .B1(new_n752_), .B2(new_n754_), .ZN(G1336gat));
  NAND4_X1  g554(.A1(new_n749_), .A2(new_n449_), .A3(new_n740_), .A4(new_n751_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G92gat), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n630_), .A2(G92gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n744_), .A2(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1337gat));
  AND2_X1   g562(.A1(new_n742_), .A2(new_n743_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n742_), .A2(new_n743_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n491_), .B(new_n444_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n744_), .A2(KEYINPUT114), .A3(new_n491_), .A4(new_n444_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n749_), .A2(new_n444_), .A3(new_n740_), .A4(new_n751_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G99gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n770_), .A2(new_n772_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1338gat));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n662_), .A2(new_n407_), .A3(new_n741_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT115), .B(new_n778_), .C1(new_n779_), .C2(new_n492_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n748_), .A2(new_n405_), .A3(new_n740_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(KEYINPUT115), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n778_), .A2(KEYINPUT115), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n781_), .A2(G106gat), .A3(new_n782_), .A4(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n744_), .A2(new_n492_), .A3(new_n405_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT53), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n780_), .A2(new_n784_), .A3(new_n788_), .A4(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n525_), .A2(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n518_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(G230gat), .A3(G233gat), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n525_), .A2(KEYINPUT117), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n791_), .B1(new_n798_), .B2(new_n535_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n535_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n804_), .B2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n531_), .A2(new_n535_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n576_), .B1(new_n802_), .B2(new_n799_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n565_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n562_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n571_), .B(new_n811_), .C1(new_n812_), .C2(new_n565_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(new_n573_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n536_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n810_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n609_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  INV_X1    g617(.A(new_n815_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n807_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n809_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n818_), .B1(new_n821_), .B2(new_n681_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n804_), .A2(new_n801_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n535_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n808_), .B(new_n814_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n826_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n614_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n817_), .A2(new_n822_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n623_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n576_), .A2(new_n489_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT116), .Z(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(new_n611_), .A3(new_n541_), .A4(new_n613_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT54), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n615_), .A2(new_n836_), .A3(new_n541_), .A4(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n405_), .B1(new_n831_), .B2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n449_), .A2(new_n447_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n444_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n278_), .B1(new_n841_), .B2(new_n576_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  INV_X1    g644(.A(new_n840_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n405_), .B(new_n846_), .C1(new_n831_), .C2(new_n838_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT59), .B1(new_n847_), .B2(new_n444_), .ZN(new_n848_));
  AND4_X1   g647(.A1(KEYINPUT59), .A2(new_n839_), .A3(new_n444_), .A4(new_n840_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n841_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n847_), .A2(KEYINPUT59), .A3(new_n444_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(KEYINPUT121), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n576_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n844_), .B1(new_n855_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g655(.A(new_n841_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n282_), .B1(new_n541_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n857_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n282_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n541_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n282_), .ZN(G1341gat));
  AOI21_X1  g660(.A(G127gat), .B1(new_n857_), .B2(new_n489_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n623_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g663(.A(G134gat), .B1(new_n857_), .B2(new_n681_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n615_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(G134gat), .ZN(G1343gat));
  AOI211_X1 g666(.A(new_n444_), .B(new_n407_), .C1(new_n831_), .C2(new_n838_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n840_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n577_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g671(.A(new_n541_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g674(.A1(new_n869_), .A2(new_n623_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT61), .B(G155gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  OAI21_X1  g677(.A(new_n594_), .B1(new_n869_), .B2(new_n609_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(KEYINPUT122), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(KEYINPUT122), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n594_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n870_), .B2(new_n882_), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n448_), .A2(new_n630_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n839_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n576_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n227_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n239_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1348gat));
  INV_X1    g690(.A(new_n885_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G176gat), .B1(new_n892_), .B2(new_n873_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n839_), .B(KEYINPUT123), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n894_), .A2(G176gat), .A3(new_n884_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n895_), .B2(new_n873_), .ZN(G1349gat));
  NOR3_X1   g695(.A1(new_n885_), .A2(new_n261_), .A3(new_n623_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n489_), .A3(new_n884_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n205_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n262_), .A3(new_n681_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G190gat), .B1(new_n885_), .B2(new_n615_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1351gat));
  NAND2_X1  g701(.A1(new_n831_), .A2(new_n838_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n412_), .A2(new_n449_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n445_), .A3(new_n904_), .ZN(new_n905_));
  OR4_X1    g704(.A1(KEYINPUT125), .A2(new_n905_), .A3(new_n247_), .A4(new_n576_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n903_), .A2(new_n445_), .A3(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n577_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n908_), .B2(new_n247_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT124), .B1(new_n908_), .B2(new_n247_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n906_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(new_n906_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n245_), .A2(KEYINPUT126), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT126), .B(G204gat), .Z(new_n915_));
  NOR2_X1   g714(.A1(new_n905_), .A2(new_n541_), .ZN(new_n916_));
  MUX2_X1   g715(.A(new_n914_), .B(new_n915_), .S(new_n916_), .Z(G1353gat));
  NOR2_X1   g716(.A1(new_n905_), .A2(new_n623_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n907_), .B2(new_n681_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n905_), .A2(new_n615_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(G218gat), .B2(new_n924_), .ZN(G1355gat));
endmodule


