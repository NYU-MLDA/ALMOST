//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n994_, new_n995_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1003_, new_n1005_,
    new_n1006_, new_n1007_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n202_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(G134gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n203_), .A2(G127gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT79), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI211_X1 g017(.A(KEYINPUT80), .B(new_n202_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT1), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n227_), .B2(KEYINPUT1), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232_));
  INV_X1    g031(.A(G155gat), .ZN(new_n233_));
  INV_X1    g032(.A(G162gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237_));
  AND2_X1   g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n235_), .A2(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n226_), .B1(new_n231_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n242_), .A2(new_n244_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n238_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n221_), .B1(new_n240_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n235_), .A2(new_n236_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT85), .B1(new_n238_), .B2(new_n237_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n238_), .A2(new_n237_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT1), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n226_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n247_), .A2(new_n248_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT86), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n220_), .A2(new_n250_), .A3(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n255_), .A2(new_n256_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n210_), .A2(new_n216_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(KEYINPUT4), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n220_), .A2(new_n250_), .A3(new_n267_), .A4(new_n259_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G85gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT0), .B(G57gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT96), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n269_), .A2(KEYINPUT96), .A3(new_n270_), .A4(new_n274_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n220_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G71gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G227gat), .A2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G15gat), .ZN(new_n288_));
  INV_X1    g087(.A(G15gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(G227gat), .A3(G233gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n290_), .A3(new_n286_), .ZN(new_n293_));
  AOI21_X1  g092(.A(G99gat), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  INV_X1    g094(.A(G99gat), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n295_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n300_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT25), .B(G183gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT26), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT75), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n311_), .A3(G190gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT74), .B1(new_n311_), .B2(G190gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n318_));
  INV_X1    g117(.A(G190gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT26), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n304_), .B(new_n309_), .C1(new_n316_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G183gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n299_), .A2(new_n301_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n325_), .C1(new_n303_), .C2(new_n299_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G169gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(KEYINPUT30), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT30), .B1(new_n322_), .B2(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n298_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n294_), .A2(new_n297_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n330_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT77), .B(G43gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n333_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n285_), .B1(new_n343_), .B2(KEYINPUT82), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n340_), .A2(new_n341_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n284_), .B2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(KEYINPUT83), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350_));
  INV_X1    g149(.A(new_n339_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n331_), .A2(new_n332_), .A3(new_n298_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n337_), .B1(new_n336_), .B2(new_n330_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n333_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT78), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n284_), .B1(new_n356_), .B2(new_n346_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n345_), .A2(new_n347_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n350_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n282_), .B1(new_n349_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n250_), .A2(new_n259_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI211_X1 g163(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n250_), .C2(new_n259_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G22gat), .B(G50gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n240_), .A2(new_n249_), .A3(new_n221_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT86), .B1(new_n257_), .B2(new_n258_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT28), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n366_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT92), .B1(new_n368_), .B2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G78gat), .B(G106gat), .Z(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT87), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G218gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G211gat), .ZN(new_n381_));
  INV_X1    g180(.A(G211gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G218gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G197gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G204gat), .ZN(new_n388_));
  INV_X1    g187(.A(G204gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G197gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n381_), .A2(new_n383_), .A3(KEYINPUT89), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n386_), .A2(KEYINPUT21), .A3(new_n391_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT21), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n381_), .A2(new_n383_), .A3(KEYINPUT89), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT89), .B1(new_n381_), .B2(new_n383_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n387_), .A3(G204gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT21), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(KEYINPUT88), .B2(new_n395_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n393_), .B(new_n394_), .C1(new_n400_), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n386_), .A2(new_n392_), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT21), .B(new_n402_), .C1(new_n391_), .C2(new_n401_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n397_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n394_), .B1(new_n409_), .B2(new_n393_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n379_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n261_), .B2(new_n363_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT90), .B(KEYINPUT29), .C1(new_n240_), .C2(new_n249_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n250_), .A2(new_n259_), .A3(KEYINPUT29), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n393_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n379_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n376_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(KEYINPUT91), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n378_), .B1(new_n422_), .B2(new_n405_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n414_), .A3(new_n413_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n376_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n420_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n367_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n372_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n375_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n426_), .A3(new_n420_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n301_), .A2(KEYINPUT76), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n301_), .A2(KEYINPUT76), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n300_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n323_), .A2(KEYINPUT25), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G183gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n319_), .A2(KEYINPUT26), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .A4(new_n312_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n309_), .A2(new_n438_), .A3(new_n325_), .A4(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n299_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n445_), .A2(new_n302_), .B1(new_n323_), .B2(new_n319_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n328_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n444_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n418_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n409_), .A2(new_n322_), .A3(new_n393_), .A4(new_n329_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(KEYINPUT20), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G226gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT19), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n334_), .B2(new_n418_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n453_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n456_), .B(new_n457_), .C1(new_n418_), .C2(new_n448_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G8gat), .B(G36gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT18), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT27), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n438_), .A2(new_n325_), .A3(new_n443_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n304_), .A2(new_n324_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n468_), .A2(new_n309_), .B1(new_n469_), .B2(new_n328_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n422_), .A2(new_n470_), .A3(new_n405_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n457_), .B1(new_n471_), .B2(new_n456_), .ZN(new_n472_));
  AND4_X1   g271(.A1(KEYINPUT20), .A2(new_n449_), .A3(new_n457_), .A4(new_n450_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT95), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n463_), .B(KEYINPUT97), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n466_), .A2(KEYINPUT27), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n467_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n435_), .A2(new_n482_), .A3(KEYINPUT98), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT98), .B1(new_n435_), .B2(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n360_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n463_), .A2(KEYINPUT32), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n459_), .B2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT32), .B(new_n463_), .C1(new_n459_), .C2(KEYINPUT94), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n477_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n282_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n269_), .A2(KEYINPUT33), .A3(new_n270_), .A4(new_n274_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n260_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n260_), .A2(KEYINPUT4), .A3(new_n263_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n268_), .A2(new_n265_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n279_), .B(new_n494_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n493_), .A2(new_n497_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n275_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n492_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n497_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n275_), .A2(new_n499_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(KEYINPUT93), .A3(new_n503_), .A4(new_n493_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n491_), .A2(new_n501_), .A3(new_n504_), .A4(new_n435_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n349_), .A2(new_n359_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n478_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n466_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n463_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI22_X1  g310(.A1(new_n508_), .A2(new_n480_), .B1(new_n511_), .B2(KEYINPUT27), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n434_), .B(new_n432_), .C1(new_n512_), .C2(new_n282_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n505_), .A2(new_n506_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n485_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G29gat), .B(G36gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT68), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(KEYINPUT68), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n519_), .A2(KEYINPUT69), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n517_), .A2(KEYINPUT68), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n523_), .B2(new_n518_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n521_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT69), .B1(new_n519_), .B2(new_n520_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n522_), .A3(new_n518_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n516_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532_));
  INV_X1    g331(.A(G1gat), .ZN(new_n533_));
  INV_X1    g332(.A(G8gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT14), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G8gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n526_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n528_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT15), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n531_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n538_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n545_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n544_), .A2(new_n538_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n515_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT10), .B(G99gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT6), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(G99gat), .B2(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT6), .ZN(new_n565_));
  OAI22_X1  g364(.A1(new_n561_), .A2(G106gat), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(G85gat), .ZN(new_n568_));
  INV_X1    g367(.A(G92gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n570_), .A2(new_n571_), .B1(new_n572_), .B2(G92gat), .ZN(new_n573_));
  AND2_X1   g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n574_), .A2(new_n575_), .A3(KEYINPUT9), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT64), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  OAI22_X1  g376(.A1(new_n574_), .A2(new_n575_), .B1(KEYINPUT9), .B2(new_n569_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT64), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n571_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n578_), .B(new_n579_), .C1(KEYINPUT9), .C2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n567_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT8), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT7), .ZN(new_n585_));
  INV_X1    g384(.A(G106gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n296_), .A3(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n584_), .B(new_n587_), .C1(new_n563_), .C2(new_n565_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT65), .B1(new_n574_), .B2(new_n575_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT65), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n570_), .A2(new_n590_), .A3(new_n571_), .ZN(new_n591_));
  AND4_X1   g390(.A1(new_n583_), .A2(new_n588_), .A3(new_n589_), .A4(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n589_), .A2(new_n591_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n583_), .B1(new_n593_), .B2(new_n588_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n582_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT11), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT11), .ZN(new_n598_));
  XOR2_X1   g397(.A(G71gat), .B(G78gat), .Z(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT12), .B1(new_n595_), .B2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n602_), .B(new_n582_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n595_), .A2(KEYINPUT66), .A3(KEYINPUT12), .A4(new_n603_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n595_), .A2(KEYINPUT12), .A3(new_n603_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT66), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n593_), .A2(new_n588_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT8), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n593_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n578_), .B1(KEYINPUT9), .B2(new_n580_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n566_), .B1(new_n618_), .B2(KEYINPUT64), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n616_), .A2(new_n617_), .B1(new_n619_), .B2(new_n581_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n602_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n614_), .B1(new_n621_), .B2(new_n606_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n613_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT67), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n613_), .A2(new_n622_), .A3(KEYINPUT67), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n613_), .A2(new_n622_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n626_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n632_), .A2(KEYINPUT13), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT13), .B1(new_n632_), .B2(new_n634_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT35), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n544_), .A2(new_n620_), .B1(new_n642_), .B2(new_n641_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT70), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n531_), .A2(new_n542_), .A3(new_n595_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n648_), .B(new_n645_), .C1(new_n646_), .C2(new_n644_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT36), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n650_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n654_), .B(KEYINPUT36), .Z(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT71), .Z(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT72), .ZN(new_n660_));
  OAI22_X1  g459(.A1(new_n656_), .A2(new_n659_), .B1(new_n660_), .B2(KEYINPUT37), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT37), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT73), .Z(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  OAI221_X1 g464(.A(new_n663_), .B1(new_n660_), .B2(KEYINPUT37), .C1(new_n656_), .C2(new_n659_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n538_), .B(new_n602_), .Z(new_n668_));
  NAND2_X1  g467(.A1(G231gat), .A2(G233gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT17), .ZN(new_n671_));
  XOR2_X1   g470(.A(G127gat), .B(G155gat), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT16), .ZN(new_n673_));
  XNOR2_X1  g472(.A(G183gat), .B(G211gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n670_), .A2(new_n671_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(KEYINPUT17), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n670_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n667_), .A2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n560_), .A2(new_n638_), .A3(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n533_), .A3(new_n282_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT38), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n637_), .A2(new_n559_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n685_), .A2(KEYINPUT99), .A3(new_n679_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT99), .B1(new_n685_), .B2(new_n679_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n688_));
  INV_X1    g487(.A(new_n659_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n650_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n656_), .A2(new_n659_), .A3(KEYINPUT100), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n485_), .B2(new_n514_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n687_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n282_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G1gat), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n684_), .A2(new_n698_), .ZN(G1324gat));
  NAND4_X1  g498(.A1(new_n686_), .A2(new_n687_), .A3(new_n695_), .A4(new_n512_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT101), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G8gat), .B1(new_n700_), .B2(KEYINPUT101), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT39), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n700_), .A2(KEYINPUT101), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT39), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(G8gat), .A4(new_n701_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n682_), .A2(new_n534_), .A3(new_n512_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(KEYINPUT40), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1325gat));
  OAI21_X1  g513(.A(G15gat), .B1(new_n696_), .B2(new_n506_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT41), .Z(new_n716_));
  INV_X1    g515(.A(new_n506_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n682_), .A2(new_n289_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1326gat));
  OAI21_X1  g518(.A(G22gat), .B1(new_n696_), .B2(new_n435_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT42), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n435_), .A2(G22gat), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT102), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n682_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1327gat));
  NOR2_X1   g524(.A1(new_n685_), .A2(new_n680_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  INV_X1    g526(.A(new_n667_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n515_), .B2(new_n728_), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT43), .B(new_n667_), .C1(new_n485_), .C2(new_n514_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(KEYINPUT103), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT103), .B1(new_n731_), .B2(new_n732_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT44), .B(new_n726_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(G29gat), .A3(new_n282_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n679_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(new_n636_), .A3(new_n635_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n515_), .A2(new_n740_), .A3(new_n559_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT104), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n515_), .A2(new_n740_), .A3(new_n743_), .A4(new_n559_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(new_n697_), .ZN(new_n746_));
  OAI22_X1  g545(.A1(new_n736_), .A2(new_n738_), .B1(G29gat), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT105), .ZN(G1328gat));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  INV_X1    g548(.A(G36gat), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n751_));
  INV_X1    g550(.A(new_n726_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n515_), .A2(new_n728_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT43), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n515_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n756_), .B2(KEYINPUT44), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n757_), .A2(new_n733_), .B1(KEYINPUT44), .B2(new_n756_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n750_), .B1(new_n758_), .B2(new_n512_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n742_), .A2(new_n750_), .A3(new_n512_), .A4(new_n744_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT106), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT106), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n761_), .A2(KEYINPUT106), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(KEYINPUT106), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(KEYINPUT45), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n749_), .B1(new_n759_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n737_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G36gat), .B1(new_n770_), .B2(new_n482_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(KEYINPUT46), .A3(new_n767_), .A4(new_n764_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(G1329gat));
  AND3_X1   g572(.A1(new_n737_), .A2(G43gat), .A3(new_n717_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n774_), .B(KEYINPUT107), .C1(new_n734_), .C2(new_n735_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT108), .B(G43gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n745_), .B2(new_n506_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT47), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n777_), .A2(new_n778_), .A3(new_n783_), .A4(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1330gat));
  INV_X1    g584(.A(G50gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n435_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n435_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n742_), .A2(new_n788_), .A3(new_n744_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n758_), .A2(new_n787_), .B1(new_n786_), .B2(new_n789_), .ZN(G1331gat));
  NOR2_X1   g589(.A1(new_n637_), .A2(new_n559_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n515_), .A2(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(new_n681_), .ZN(new_n793_));
  AOI211_X1 g592(.A(G57gat), .B(new_n697_), .C1(new_n793_), .C2(KEYINPUT109), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(KEYINPUT109), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n680_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(new_n282_), .A3(new_n695_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n794_), .A2(new_n795_), .B1(G57gat), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT110), .ZN(G1332gat));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n695_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G64gat), .B1(new_n801_), .B2(new_n482_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT48), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n482_), .A2(G64gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n793_), .B2(new_n804_), .ZN(G1333gat));
  OAI21_X1  g604(.A(G71gat), .B1(new_n801_), .B2(new_n506_), .ZN(new_n806_));
  XOR2_X1   g605(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n717_), .A2(new_n286_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n793_), .B2(new_n809_), .ZN(G1334gat));
  OAI21_X1  g609(.A(G78gat), .B1(new_n801_), .B2(new_n435_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT50), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n435_), .A2(G78gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n793_), .B2(new_n813_), .ZN(G1335gat));
  NOR2_X1   g613(.A1(new_n792_), .A2(new_n739_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n568_), .A3(new_n282_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n754_), .A2(new_n817_), .A3(new_n755_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT112), .B1(new_n729_), .B2(new_n730_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n559_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n679_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT113), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n818_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n282_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n816_), .B1(new_n824_), .B2(new_n568_), .ZN(G1336gat));
  NAND3_X1  g624(.A1(new_n815_), .A2(new_n569_), .A3(new_n512_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n823_), .A2(new_n512_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n569_), .ZN(G1337gat));
  NOR2_X1   g627(.A1(new_n506_), .A2(new_n561_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n815_), .A2(new_n829_), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT115), .Z(new_n831_));
  NAND4_X1  g630(.A1(new_n818_), .A2(new_n819_), .A3(new_n717_), .A4(new_n822_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G99gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G99gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n837_));
  OR2_X1    g636(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n832_), .A2(G99gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT114), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n832_), .A2(new_n833_), .A3(G99gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(KEYINPUT116), .A3(KEYINPUT51), .A4(new_n831_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n839_), .A2(new_n844_), .ZN(G1338gat));
  NAND3_X1  g644(.A1(new_n815_), .A2(new_n586_), .A3(new_n788_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n729_), .A2(new_n730_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n822_), .A2(new_n788_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G106gat), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT117), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n852_), .B(G106gat), .C1(new_n847_), .C2(new_n848_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n851_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n846_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT53), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n858_), .B(new_n846_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1339gat));
  OR2_X1    g659(.A1(new_n483_), .A2(new_n484_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n282_), .A3(new_n717_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n632_), .A2(new_n559_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT12), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n620_), .B2(new_n602_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n612_), .A2(new_n605_), .A3(new_n609_), .A4(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n614_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT55), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n613_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n869_), .A2(new_n873_), .A3(new_n614_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT56), .B1(new_n876_), .B2(new_n626_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n869_), .B2(new_n614_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n613_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT56), .B(new_n626_), .C1(new_n880_), .C2(new_n874_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n866_), .B1(new_n877_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n632_), .A2(new_n634_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n549_), .A2(new_n550_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n556_), .B1(new_n886_), .B2(new_n548_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n543_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n887_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(KEYINPUT118), .A3(new_n888_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n884_), .A2(new_n558_), .A3(new_n890_), .A4(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n883_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894_), .B2(new_n693_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n626_), .B1(new_n880_), .B2(new_n874_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n865_), .B1(new_n898_), .B2(new_n881_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n890_), .A3(new_n558_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n634_), .B2(new_n632_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n693_), .C1(new_n899_), .C2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n895_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n876_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n626_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n881_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n907_), .A3(new_n898_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n900_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n908_), .A2(KEYINPUT58), .A3(new_n909_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n728_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n680_), .B1(new_n904_), .B2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n637_), .A2(new_n667_), .A3(new_n820_), .A4(new_n680_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT54), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n863_), .B(new_n864_), .C1(new_n914_), .C2(new_n917_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n908_), .A2(KEYINPUT58), .A3(new_n909_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n919_), .A2(new_n910_), .A3(new_n667_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n693_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n902_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n679_), .B1(new_n920_), .B2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n862_), .B1(new_n925_), .B2(new_n916_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n927_));
  OAI21_X1  g726(.A(new_n918_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G113gat), .B1(new_n928_), .B2(new_n820_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n926_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n820_), .A2(G113gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1340gat));
  NOR2_X1   g731(.A1(new_n637_), .A2(KEYINPUT60), .ZN(new_n933_));
  MUX2_X1   g732(.A(new_n933_), .B(KEYINPUT60), .S(G120gat), .Z(new_n934_));
  NAND2_X1  g733(.A1(new_n926_), .A2(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT121), .ZN(new_n936_));
  OAI21_X1  g735(.A(G120gat), .B1(new_n928_), .B2(new_n637_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1341gat));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939_));
  AOI211_X1 g738(.A(new_n679_), .B(new_n862_), .C1(new_n925_), .C2(new_n916_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(G127gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n679_), .A2(new_n205_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n918_), .B(new_n942_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n925_), .A2(new_n916_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n944_), .A2(new_n680_), .A3(new_n863_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n945_), .A2(KEYINPUT122), .A3(new_n205_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n941_), .A2(new_n943_), .A3(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n941_), .A2(new_n943_), .A3(new_n946_), .A4(KEYINPUT123), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1342gat));
  OAI21_X1  g750(.A(G134gat), .B1(new_n928_), .B2(new_n667_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n926_), .A2(new_n203_), .A3(new_n694_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1343gat));
  NOR2_X1   g753(.A1(new_n717_), .A2(new_n435_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n956_), .B1(new_n925_), .B2(new_n916_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n697_), .A2(new_n512_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n820_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(new_n222_), .ZN(G1344gat));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n637_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(new_n223_), .ZN(G1345gat));
  NOR2_X1   g762(.A1(new_n959_), .A2(new_n679_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT61), .B(G155gat), .ZN(new_n965_));
  XOR2_X1   g764(.A(new_n964_), .B(new_n965_), .Z(G1346gat));
  NOR3_X1   g765(.A1(new_n959_), .A2(new_n234_), .A3(new_n667_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n957_), .A2(new_n694_), .A3(new_n958_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n234_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n968_), .A2(KEYINPUT124), .A3(new_n234_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n967_), .B1(new_n971_), .B2(new_n972_), .ZN(G1347gat));
  NOR2_X1   g772(.A1(new_n482_), .A2(new_n282_), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n975_), .A2(new_n506_), .ZN(new_n976_));
  NAND4_X1  g775(.A1(new_n944_), .A2(new_n559_), .A3(new_n435_), .A4(new_n976_), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978_));
  AND3_X1   g777(.A1(new_n977_), .A2(new_n978_), .A3(G169gat), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n977_), .B2(G169gat), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n944_), .A2(new_n435_), .A3(new_n976_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(KEYINPUT22), .B(G169gat), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n559_), .A2(new_n982_), .ZN(new_n983_));
  XOR2_X1   g782(.A(new_n983_), .B(KEYINPUT125), .Z(new_n984_));
  OAI22_X1  g783(.A1(new_n979_), .A2(new_n980_), .B1(new_n981_), .B2(new_n984_), .ZN(G1348gat));
  NAND2_X1  g784(.A1(new_n944_), .A2(new_n435_), .ZN(new_n986_));
  OR2_X1    g785(.A1(new_n986_), .A2(KEYINPUT126), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(KEYINPUT126), .ZN(new_n988_));
  INV_X1    g787(.A(G176gat), .ZN(new_n989_));
  NOR4_X1   g788(.A1(new_n637_), .A2(new_n989_), .A3(new_n506_), .A4(new_n975_), .ZN(new_n990_));
  NAND3_X1  g789(.A1(new_n987_), .A2(new_n988_), .A3(new_n990_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n989_), .B1(new_n981_), .B2(new_n637_), .ZN(new_n992_));
  AND2_X1   g791(.A1(new_n991_), .A2(new_n992_), .ZN(G1349gat));
  NOR3_X1   g792(.A1(new_n981_), .A2(new_n679_), .A3(new_n310_), .ZN(new_n994_));
  NAND4_X1  g793(.A1(new_n987_), .A2(new_n680_), .A3(new_n976_), .A4(new_n988_), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n994_), .B1(new_n995_), .B2(new_n323_), .ZN(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n981_), .B2(new_n667_), .ZN(new_n997_));
  NAND3_X1  g796(.A1(new_n694_), .A2(new_n442_), .A3(new_n312_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n997_), .B1(new_n981_), .B2(new_n998_), .ZN(G1351gat));
  AOI211_X1 g798(.A(new_n956_), .B(new_n975_), .C1(new_n925_), .C2(new_n916_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n1000_), .A2(new_n559_), .ZN(new_n1001_));
  XNOR2_X1  g800(.A(new_n1001_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g801(.A1(new_n1000_), .A2(new_n638_), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(new_n1003_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g803(.A1(new_n1000_), .A2(new_n680_), .ZN(new_n1005_));
  OAI21_X1  g804(.A(new_n1005_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1006_));
  XOR2_X1   g805(.A(KEYINPUT63), .B(G211gat), .Z(new_n1007_));
  OAI21_X1  g806(.A(new_n1006_), .B1(new_n1005_), .B2(new_n1007_), .ZN(G1354gat));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009_));
  NOR2_X1   g808(.A1(new_n693_), .A2(G218gat), .ZN(new_n1010_));
  NAND2_X1  g809(.A1(new_n1000_), .A2(new_n1010_), .ZN(new_n1011_));
  AND2_X1   g810(.A1(new_n1000_), .A2(new_n728_), .ZN(new_n1012_));
  OAI211_X1 g811(.A(new_n1009_), .B(new_n1011_), .C1(new_n1012_), .C2(new_n380_), .ZN(new_n1013_));
  INV_X1    g812(.A(new_n1011_), .ZN(new_n1014_));
  AOI21_X1  g813(.A(new_n380_), .B1(new_n1000_), .B2(new_n728_), .ZN(new_n1015_));
  OAI21_X1  g814(.A(KEYINPUT127), .B1(new_n1014_), .B2(new_n1015_), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1013_), .A2(new_n1016_), .ZN(G1355gat));
endmodule


