//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT86), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT87), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT87), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G155gat), .A3(G162gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT88), .B1(new_n208_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n211_), .A2(new_n213_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n207_), .B(new_n216_), .C1(new_n217_), .C2(new_n209_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n209_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G141gat), .ZN(new_n221_));
  INV_X1    g020(.A(G148gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(KEYINPUT2), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .A4(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n217_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n207_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237_));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n235_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT97), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(KEYINPUT97), .A3(new_n243_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(KEYINPUT4), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n240_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G85gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n258_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n252_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G8gat), .B(G36gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(G197gat), .A2(G204gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G218gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(G211gat), .ZN(new_n278_));
  INV_X1    g077(.A(G211gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT91), .B1(new_n279_), .B2(G218gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n276_), .B(KEYINPUT21), .C1(new_n278_), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(KEYINPUT21), .A3(new_n274_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n280_), .A2(new_n278_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT23), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(G183gat), .B2(G190gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT84), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n290_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  INV_X1    g104(.A(G176gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(KEYINPUT82), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT82), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(G169gat), .B2(G176gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT24), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n293_), .A2(new_n295_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT25), .B(G183gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT26), .B(G190gat), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI211_X1 g113(.A(new_n310_), .B(new_n311_), .C1(new_n312_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n307_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(G169gat), .B2(G176gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n288_), .B1(new_n304_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT81), .B(G190gat), .Z(new_n325_));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n312_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n320_), .B1(new_n330_), .B2(new_n317_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n297_), .A2(new_n299_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n293_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n329_), .A2(new_n322_), .A3(new_n331_), .A4(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n325_), .A2(new_n291_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n290_), .B1(new_n336_), .B2(new_n311_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n281_), .A2(new_n286_), .A3(KEYINPUT92), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT92), .B1(new_n281_), .B2(new_n286_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n324_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT99), .B(KEYINPUT20), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n287_), .B1(new_n315_), .B2(new_n322_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n302_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n338_), .A2(new_n341_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n272_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT100), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(KEYINPUT100), .B(new_n272_), .C1(new_n347_), .C2(new_n352_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n346_), .B1(new_n324_), .B2(new_n342_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n304_), .A2(new_n288_), .A3(new_n323_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n358_), .A2(new_n351_), .A3(KEYINPUT20), .A4(new_n345_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n355_), .A2(new_n356_), .B1(new_n360_), .B2(new_n271_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n265_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT101), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n263_), .A2(new_n262_), .A3(new_n259_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT33), .B1(new_n365_), .B2(KEYINPUT98), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n270_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n357_), .A2(new_n270_), .A3(new_n359_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n251_), .A2(new_n252_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n246_), .A2(new_n247_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n258_), .B1(new_n370_), .B2(new_n253_), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n367_), .B(new_n368_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT98), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT33), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n261_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n265_), .A2(new_n361_), .A3(KEYINPUT101), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n364_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT93), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT28), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n242_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n242_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G22gat), .B(G50gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n386_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n389_), .B1(new_n390_), .B2(new_n384_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n341_), .B1(new_n242_), .B2(new_n383_), .ZN(new_n392_));
  INV_X1    g191(.A(G228gat), .ZN(new_n393_));
  INV_X1    g192(.A(G233gat), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n394_), .A2(KEYINPUT89), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(KEYINPUT89), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT90), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n288_), .A2(new_n398_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n242_), .B2(new_n383_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n388_), .A2(new_n391_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n381_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n391_), .A2(new_n388_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n380_), .A3(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n378_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n270_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n357_), .A2(new_n270_), .A3(new_n359_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(KEYINPUT27), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT102), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT27), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n368_), .B2(new_n367_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT102), .A4(KEYINPUT27), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n410_), .A2(new_n265_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n411_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426_));
  INV_X1    g225(.A(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT30), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n338_), .B(new_n429_), .Z(new_n430_));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(G15gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n338_), .B(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n433_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(KEYINPUT85), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT31), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT31), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n435_), .A2(KEYINPUT85), .A3(new_n440_), .A4(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n243_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n239_), .A3(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT103), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n406_), .A2(new_n409_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n421_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n265_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n419_), .A2(new_n420_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(new_n410_), .A3(KEYINPUT103), .A4(new_n417_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT104), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n445_), .B1(new_n456_), .B2(new_n446_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n457_), .A2(KEYINPUT104), .A3(new_n450_), .A4(new_n452_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n425_), .A2(new_n445_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G29gat), .B(G36gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n460_), .A2(new_n461_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G43gat), .B(G50gat), .Z(new_n464_));
  OR3_X1    g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT80), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT77), .B(G1gat), .ZN(new_n469_));
  INV_X1    g268(.A(G8gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT14), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G1gat), .B(G8gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n468_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n467_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n465_), .A2(KEYINPUT15), .A3(new_n466_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(new_n475_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n468_), .A2(new_n475_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n477_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n479_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G141gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n479_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n459_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT13), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G85gat), .B(G92gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT6), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n499_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT67), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n499_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n505_), .A2(new_n507_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514_));
  INV_X1    g313(.A(G99gat), .ZN(new_n515_));
  INV_X1    g314(.A(G106gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n500_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n512_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT8), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n503_), .A2(KEYINPUT65), .A3(new_n508_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n499_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n511_), .A2(new_n521_), .A3(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT64), .B(G85gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G92gat), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n530_), .A2(KEYINPUT9), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n512_), .A2(KEYINPUT9), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT10), .B(G99gat), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n516_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n532_), .A2(new_n533_), .A3(new_n535_), .A4(new_n508_), .ZN(new_n536_));
  OR2_X1    g335(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G78gat), .ZN(new_n540_));
  INV_X1    g339(.A(G78gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n541_), .A3(new_n538_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n540_), .A2(new_n542_), .B1(KEYINPUT11), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(KEYINPUT11), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n540_), .A2(new_n542_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n528_), .A2(new_n536_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT70), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n528_), .A2(new_n536_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n547_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n553_), .A2(new_n554_), .B1(KEYINPUT70), .B2(new_n549_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(KEYINPUT70), .ZN(new_n556_));
  AOI211_X1 g355(.A(new_n556_), .B(new_n547_), .C1(new_n528_), .C2(new_n536_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n551_), .B(new_n552_), .C1(new_n555_), .C2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n547_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n548_), .A2(KEYINPUT69), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n558_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n558_), .A2(new_n563_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n567_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(KEYINPUT72), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT72), .B1(new_n571_), .B2(new_n573_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n498_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n574_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n553_), .A2(new_n467_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n483_), .A2(new_n553_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n481_), .A2(new_n482_), .B1(new_n536_), .B2(new_n528_), .ZN(new_n589_));
  OAI211_X1 g388(.A(KEYINPUT35), .B(new_n585_), .C1(new_n581_), .C2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n590_), .A3(KEYINPUT75), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT74), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n588_), .A2(new_n590_), .A3(KEYINPUT75), .A4(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n588_), .A2(new_n590_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n598_), .A2(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT76), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT76), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n602_), .A2(KEYINPUT76), .A3(new_n603_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n475_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n554_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT79), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n612_), .A2(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n619_), .A3(new_n612_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n580_), .A2(new_n609_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n497_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n469_), .A3(new_n265_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  INV_X1    g427(.A(new_n602_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n459_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n623_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n577_), .A2(new_n579_), .A3(new_n495_), .A4(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT106), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n265_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n627_), .A2(new_n628_), .B1(new_n636_), .B2(G1gat), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n627_), .A2(new_n628_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT105), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(KEYINPUT105), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(G1324gat));
  NAND3_X1  g440(.A1(new_n630_), .A2(new_n633_), .A3(new_n421_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT107), .B1(new_n642_), .B2(G8gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n642_), .A2(G8gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n644_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n421_), .A2(new_n470_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n625_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n648_), .A2(KEYINPUT40), .A3(new_n649_), .A4(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n647_), .A2(new_n646_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n649_), .A2(new_n651_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n657_), .ZN(G1325gat));
  NAND2_X1  g457(.A1(new_n635_), .A2(new_n449_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G15gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT108), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n662_), .A3(G15gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(KEYINPUT41), .A3(new_n663_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n626_), .A2(new_n432_), .A3(new_n449_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(G1326gat));
  OR3_X1    g468(.A1(new_n625_), .A2(G22gat), .A3(new_n410_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G22gat), .B1(new_n634_), .B2(new_n410_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(KEYINPUT42), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(KEYINPUT42), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT109), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n670_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n629_), .A2(new_n623_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n580_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n497_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n265_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n608_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n685_), .B2(KEYINPUT110), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n459_), .B2(new_n685_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n455_), .A2(new_n458_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n378_), .A2(new_n410_), .B1(new_n423_), .B2(new_n422_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n449_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n609_), .B(new_n686_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n580_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n495_), .A3(new_n623_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n698_), .B(new_n695_), .C1(new_n688_), .C2(new_n692_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n265_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n682_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n700_), .B2(new_n421_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n497_), .A2(new_n704_), .A3(new_n421_), .A4(new_n680_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n705_), .B2(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n697_), .A2(new_n699_), .A3(new_n422_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT46), .B(new_n707_), .C1(new_n710_), .C2(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1329gat));
  NOR4_X1   g511(.A1(new_n697_), .A2(new_n699_), .A3(new_n427_), .A4(new_n445_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G43gat), .B1(new_n681_), .B2(new_n449_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT47), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n445_), .A2(new_n427_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n700_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n719_), .ZN(G1330gat));
  AOI21_X1  g519(.A(G50gat), .B1(new_n681_), .B2(new_n447_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n447_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n700_), .B2(new_n722_), .ZN(G1331gat));
  NOR3_X1   g522(.A1(new_n694_), .A2(new_n495_), .A3(new_n623_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n630_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(G57gat), .A3(new_n265_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n459_), .A2(new_n495_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n609_), .A2(new_n623_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n580_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT111), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n265_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n734_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n727_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n738_), .A3(new_n421_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n726_), .A2(new_n421_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(G64gat), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G64gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n725_), .B2(new_n445_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT49), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n445_), .A2(G71gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT114), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n732_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1334gat));
  NAND3_X1  g549(.A1(new_n732_), .A2(new_n541_), .A3(new_n447_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G78gat), .B1(new_n725_), .B2(new_n410_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT50), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT50), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT115), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n751_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n694_), .A2(new_n679_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n728_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n265_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n688_), .A2(new_n692_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n694_), .A2(new_n495_), .A3(new_n631_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n450_), .A2(new_n530_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n762_), .B1(new_n766_), .B2(new_n767_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n531_), .A3(new_n421_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n763_), .A2(new_n422_), .A3(new_n765_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n531_), .ZN(G1337gat));
  AOI21_X1  g570(.A(new_n515_), .B1(new_n766_), .B2(new_n449_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n728_), .A2(new_n449_), .A3(new_n534_), .A4(new_n760_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT116), .ZN(new_n774_));
  OR3_X1    g573(.A1(new_n772_), .A2(KEYINPUT51), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n772_), .B2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n761_), .A2(new_n516_), .A3(new_n447_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n693_), .A2(new_n447_), .A3(new_n764_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n516_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n786_), .B(new_n778_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n495_), .A2(new_n571_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n551_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n552_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(KEYINPUT55), .A3(new_n558_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n555_), .A2(new_n557_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n552_), .A4(new_n551_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n794_), .A2(KEYINPUT119), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT119), .B1(new_n794_), .B2(new_n797_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n567_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT56), .B(new_n567_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n790_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n476_), .A2(new_n477_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n485_), .A2(new_n486_), .A3(new_n478_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n492_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n494_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n578_), .B2(new_n574_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n602_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n808_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n571_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n685_), .B1(new_n813_), .B2(KEYINPUT58), .ZN(new_n814_));
  INV_X1    g613(.A(new_n812_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n794_), .A2(new_n797_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n794_), .A2(KEYINPUT119), .A3(new_n797_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n567_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n803_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n815_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n789_), .A2(new_n810_), .B1(new_n814_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n790_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n811_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n629_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT57), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n631_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n729_), .A2(new_n496_), .A3(new_n577_), .A4(new_n579_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n832_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n457_), .A2(new_n265_), .A3(new_n452_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT58), .B(new_n815_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n609_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n813_), .A2(KEYINPUT58), .ZN(new_n846_));
  OAI22_X1  g645(.A1(new_n830_), .A2(KEYINPUT57), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n814_), .A2(new_n825_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(KEYINPUT120), .C1(KEYINPUT57), .C2(new_n830_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n831_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n839_), .B1(new_n852_), .B2(new_n623_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n842_), .A2(new_n843_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n496_), .ZN(new_n856_));
  INV_X1    g655(.A(G113gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n842_), .A2(new_n857_), .A3(new_n495_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1340gat));
  OAI21_X1  g658(.A(G120gat), .B1(new_n855_), .B2(new_n694_), .ZN(new_n860_));
  INV_X1    g659(.A(G120gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n694_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n842_), .B(new_n862_), .C1(KEYINPUT60), .C2(new_n861_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n855_), .B2(new_n623_), .ZN(new_n865_));
  INV_X1    g664(.A(G127gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n842_), .A2(new_n866_), .A3(new_n631_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1342gat));
  OAI21_X1  g667(.A(G134gat), .B1(new_n855_), .B2(new_n685_), .ZN(new_n869_));
  INV_X1    g668(.A(G134gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n842_), .A2(new_n870_), .A3(new_n629_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1343gat));
  OR2_X1    g671(.A1(new_n832_), .A2(new_n839_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n449_), .A2(new_n450_), .A3(new_n410_), .A4(new_n421_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n495_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n580_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n631_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  NOR2_X1   g681(.A1(new_n602_), .A2(G162gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n875_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n873_), .A2(new_n609_), .A3(new_n874_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n203_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT121), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n884_), .B(new_n889_), .C1(new_n886_), .C2(new_n203_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1347gat));
  NOR3_X1   g690(.A1(new_n422_), .A2(new_n445_), .A3(new_n265_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n495_), .ZN(new_n893_));
  AND2_X1   g692(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OR4_X1    g695(.A1(new_n447_), .A2(new_n853_), .A3(new_n893_), .A4(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n893_), .A2(KEYINPUT122), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n893_), .A2(KEYINPUT122), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n410_), .A3(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n831_), .B1(new_n826_), .B2(KEYINPUT120), .ZN(new_n902_));
  INV_X1    g701(.A(new_n851_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n623_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n839_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n901_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n305_), .B1(new_n906_), .B2(KEYINPUT123), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n853_), .B2(new_n901_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n898_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n901_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n847_), .A2(new_n848_), .B1(KEYINPUT57), .B2(new_n830_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n631_), .B1(new_n912_), .B2(new_n851_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT123), .B(new_n911_), .C1(new_n913_), .C2(new_n839_), .ZN(new_n914_));
  AND4_X1   g713(.A1(new_n898_), .A2(new_n909_), .A3(G169gat), .A4(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n897_), .B1(new_n910_), .B2(new_n915_), .ZN(G1348gat));
  NAND3_X1  g715(.A1(new_n580_), .A2(G176gat), .A3(new_n892_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n840_), .A2(new_n447_), .A3(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n410_), .B(new_n892_), .C1(new_n913_), .C2(new_n839_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n306_), .B1(new_n919_), .B2(new_n694_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT124), .B(new_n306_), .C1(new_n919_), .C2(new_n694_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n918_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  NAND4_X1  g723(.A1(new_n873_), .A2(new_n410_), .A3(new_n631_), .A4(new_n892_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n291_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n623_), .A2(new_n312_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n919_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n926_), .B(KEYINPUT125), .C1(new_n919_), .C2(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n919_), .B2(new_n685_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n629_), .A2(new_n314_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n919_), .B2(new_n934_), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n423_), .A2(new_n445_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n422_), .B1(new_n937_), .B2(KEYINPUT126), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n938_), .B1(KEYINPUT126), .B2(new_n937_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n840_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n495_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n580_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n631_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n945_), .A2(new_n946_), .A3(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  NAND3_X1  g748(.A1(new_n940_), .A2(new_n277_), .A3(new_n629_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n840_), .A2(new_n685_), .A3(new_n939_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n277_), .ZN(G1355gat));
endmodule


