//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G8gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G226gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT19), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT81), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT22), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G169gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n214_), .B1(new_n217_), .B2(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n213_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(G176gat), .B1(new_n216_), .B2(new_n214_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n224_), .B(KEYINPUT82), .C1(new_n214_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n227_), .B(KEYINPUT79), .Z(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT23), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT23), .B1(new_n232_), .B2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(G183gat), .B2(G190gat), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n223_), .A2(new_n226_), .A3(KEYINPUT83), .A4(new_n228_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n231_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n235_), .B(KEYINPUT80), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n234_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n215_), .A2(new_n221_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT24), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT26), .B(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT78), .B1(new_n245_), .B2(G183gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT25), .B(G183gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n244_), .B(new_n246_), .C1(new_n247_), .C2(KEYINPUT78), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n242_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n241_), .A2(new_n243_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n239_), .A2(KEYINPUT84), .A3(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G211gat), .B(G218gat), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT90), .B1(new_n258_), .B2(G197gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(G204gat), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n259_), .A2(new_n262_), .B1(G197gat), .B2(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n257_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n256_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n261_), .B2(G204gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n258_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(G204gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT21), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT91), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n262_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n258_), .A2(G197gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n264_), .A3(new_n275_), .ZN(new_n276_));
  AND4_X1   g075(.A1(KEYINPUT91), .A2(new_n276_), .A3(new_n272_), .A4(new_n257_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n265_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT94), .B1(new_n255_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n239_), .A2(KEYINPUT84), .A3(new_n250_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT84), .B1(new_n239_), .B2(new_n250_), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT94), .B(new_n278_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n241_), .B1(G183gat), .B2(G190gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n225_), .A2(new_n221_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n241_), .B(KEYINPUT93), .C1(G183gat), .C2(G190gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .A4(new_n228_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n242_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n247_), .A2(new_n244_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n236_), .A2(new_n291_), .A3(new_n243_), .A4(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT20), .B1(new_n294_), .B2(new_n278_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n212_), .B1(new_n284_), .B2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n280_), .A2(new_n281_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n276_), .A2(new_n272_), .A3(new_n257_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT91), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n266_), .A2(KEYINPUT91), .A3(new_n272_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n302_), .A3(new_n265_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n294_), .A2(new_n278_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(KEYINPUT20), .A4(new_n211_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n209_), .B1(new_n296_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT94), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n295_), .B1(new_n309_), .B2(new_n282_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n209_), .B(new_n305_), .C1(new_n310_), .C2(new_n211_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n203_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G85gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT0), .ZN(new_n316_));
  INV_X1    g115(.A(G57gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(G155gat), .B(G162gat), .Z(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(KEYINPUT86), .B2(KEYINPUT3), .ZN(new_n323_));
  INV_X1    g122(.A(G141gat), .ZN(new_n324_));
  INV_X1    g123(.A(G148gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n322_), .A2(KEYINPUT3), .ZN(new_n327_));
  OAI221_X1 g126(.A(new_n322_), .B1(KEYINPUT86), .B2(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n330_), .B(KEYINPUT2), .Z(new_n331_));
  OAI21_X1  g130(.A(new_n321_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G155gat), .ZN(new_n333_));
  INV_X1    g132(.A(G162gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT1), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(G155gat), .A3(G162gat), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n335_), .B(new_n337_), .C1(G155gat), .C2(G162gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n324_), .A2(new_n325_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n330_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n332_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342_));
  INV_X1    g141(.A(G113gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G113gat), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n344_), .A2(G120gat), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(G120gat), .B1(new_n344_), .B2(new_n346_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT96), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n341_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n347_), .A2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n332_), .A2(new_n340_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT4), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(KEYINPUT96), .A3(new_n353_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n320_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n349_), .B(new_n353_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n320_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n319_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n320_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n341_), .A2(new_n349_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n356_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n351_), .A2(KEYINPUT4), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n361_), .A3(new_n318_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n363_), .A2(KEYINPUT98), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT98), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n368_), .A2(new_n371_), .A3(new_n318_), .A4(new_n361_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n305_), .B1(new_n310_), .B2(new_n211_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n208_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n303_), .A2(new_n304_), .A3(KEYINPUT20), .A4(new_n212_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n310_), .B2(new_n212_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n209_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n379_), .A3(KEYINPUT27), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n313_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n302_), .B2(new_n265_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AND4_X1   g185(.A1(KEYINPUT88), .A2(new_n278_), .A3(new_n382_), .A4(new_n385_), .ZN(new_n387_));
  OAI21_X1  g186(.A(G78gat), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n278_), .A2(KEYINPUT88), .A3(new_n385_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(G228gat), .A3(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(G78gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n388_), .A2(G106gat), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(G106gat), .B1(new_n388_), .B2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT92), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n393_), .ZN(new_n397_));
  INV_X1    g196(.A(G106gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n388_), .A2(new_n393_), .A3(G106gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n403_));
  INV_X1    g202(.A(G50gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT28), .B(G22gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n396_), .A2(new_n402_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n399_), .A2(new_n409_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT31), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n297_), .A2(new_n349_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n255_), .A2(new_n352_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n297_), .A2(new_n349_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n255_), .A2(new_n352_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G71gat), .B(G99gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n417_), .A2(new_n426_), .A3(new_n421_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n381_), .A2(new_n412_), .A3(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n381_), .A2(new_n412_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n318_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT97), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n320_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(KEYINPUT97), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n369_), .B(KEYINPUT33), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n376_), .A2(new_n311_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n208_), .A2(KEYINPUT32), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n378_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n375_), .A2(new_n440_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n373_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n444_), .A3(new_n411_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n428_), .A2(KEYINPUT85), .A3(new_n429_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT85), .B1(new_n428_), .B2(new_n429_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT99), .B1(new_n432_), .B2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n445_), .A2(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n381_), .A2(new_n412_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT99), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n431_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G190gat), .B(G218gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT72), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G134gat), .B(G162gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT10), .B(G99gat), .Z(new_n463_));
  AND2_X1   g262(.A1(new_n463_), .A2(new_n398_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(KEYINPUT6), .Z(new_n466_));
  INV_X1    g265(.A(G85gat), .ZN(new_n467_));
  INV_X1    g266(.A(G92gat), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT9), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n464_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G85gat), .B(G92gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT9), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT64), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n474_), .B(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT65), .B(new_n471_), .C1(new_n477_), .C2(new_n466_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT8), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT67), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n473_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G43gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G50gat), .ZN(new_n488_));
  INV_X1    g287(.A(G43gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n486_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n404_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT15), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n491_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT15), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n483_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT70), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n493_), .A2(new_n479_), .A3(new_n473_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n500_), .A2(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n505_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n496_), .A2(new_n507_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n460_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n459_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n462_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT73), .B1(new_n506_), .B2(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(new_n462_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n455_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT66), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G71gat), .B(G78gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n524_));
  INV_X1    g323(.A(new_n522_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(KEYINPUT11), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n483_), .A2(new_n529_), .A3(KEYINPUT12), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n479_), .A2(new_n473_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n527_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n527_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n531_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G176gat), .B(G204gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n541_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT13), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552_));
  INV_X1    g351(.A(G8gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G1gat), .B(G8gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n495_), .A2(new_n558_), .A3(new_n492_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n493_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT75), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n493_), .B(new_n557_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT77), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n215_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G197gat), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT76), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n566_), .B(new_n569_), .C1(new_n575_), .C2(new_n574_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n551_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n557_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(new_n527_), .Z(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n232_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G211gat), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n528_), .A3(KEYINPUT17), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(KEYINPUT17), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n583_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n580_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT100), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(KEYINPUT100), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n518_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n202_), .B1(new_n597_), .B2(new_n373_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT101), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT37), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(KEYINPUT37), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n516_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n513_), .A2(new_n515_), .A3(new_n600_), .A4(KEYINPUT37), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n603_), .A2(new_n593_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n580_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n455_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n202_), .A3(new_n373_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT38), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n599_), .A2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n518_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n313_), .A2(new_n380_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n618_), .B(G8gat), .C1(new_n613_), .C2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n608_), .A2(new_n553_), .A3(new_n614_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n612_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(KEYINPUT40), .A3(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1325gat));
  INV_X1    g428(.A(G15gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n448_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n597_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n608_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n613_), .B2(new_n411_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  INV_X1    g438(.A(G22gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n608_), .A2(new_n640_), .A3(new_n412_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT104), .ZN(G1327gat));
  NOR2_X1   g442(.A1(new_n516_), .A2(new_n593_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n455_), .A2(new_n607_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n373_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n603_), .A2(new_n604_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n431_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n451_), .A2(new_n453_), .A3(new_n452_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n453_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n648_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n607_), .A2(new_n593_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n455_), .A2(KEYINPUT43), .A3(new_n649_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n655_), .B1(new_n654_), .B2(new_n648_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT44), .B(new_n658_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n660_), .A2(G29gat), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n647_), .B1(new_n664_), .B2(new_n373_), .ZN(G1328gat));
  NOR2_X1   g464(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT107), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n614_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G36gat), .B1(new_n668_), .B2(new_n659_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT105), .B(G36gat), .C1(new_n668_), .C2(new_n659_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n646_), .A2(new_n674_), .A3(new_n614_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n667_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n667_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n676_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n678_), .B(new_n679_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n677_), .A2(new_n680_), .ZN(G1329gat));
  INV_X1    g480(.A(new_n430_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n660_), .A2(G43gat), .A3(new_n682_), .A4(new_n663_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G43gat), .B1(new_n646_), .B2(new_n631_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n646_), .B2(new_n412_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n660_), .A2(G50gat), .A3(new_n663_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n412_), .ZN(G1331gat));
  INV_X1    g489(.A(new_n551_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n579_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n654_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n606_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n373_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n317_), .A2(KEYINPUT108), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n518_), .A2(new_n593_), .A3(new_n693_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n317_), .B1(new_n373_), .B2(KEYINPUT108), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n697_), .B2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n698_), .B2(new_n615_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT48), .Z(new_n703_));
  INV_X1    g502(.A(new_n695_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(G64gat), .A3(new_n615_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n698_), .B2(new_n448_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT49), .Z(new_n708_));
  NOR3_X1   g507(.A1(new_n704_), .A2(G71gat), .A3(new_n448_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1334gat));
  OAI21_X1  g509(.A(G78gat), .B1(new_n698_), .B2(new_n411_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT50), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n411_), .A2(G78gat), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT109), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n704_), .B2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n694_), .A2(new_n645_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n373_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT110), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n657_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n593_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n693_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n650_), .A2(KEYINPUT111), .A3(new_n656_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n373_), .A2(G85gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n718_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1336gat));
  NOR3_X1   g528(.A1(new_n725_), .A2(new_n468_), .A3(new_n615_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G92gat), .B1(new_n716_), .B2(new_n614_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1337gat));
  NAND3_X1  g531(.A1(new_n716_), .A2(new_n463_), .A3(new_n682_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT113), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n720_), .A2(new_n631_), .A3(new_n723_), .A4(new_n724_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G99gat), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n737_));
  AND3_X1   g536(.A1(new_n734_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT115), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT115), .B1(new_n738_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1338gat));
  AOI211_X1 g542(.A(new_n411_), .B(new_n722_), .C1(new_n650_), .C2(new_n656_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT116), .B1(new_n744_), .B2(new_n398_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n657_), .A2(new_n412_), .A3(new_n723_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT52), .A3(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n716_), .A2(new_n398_), .A3(new_n412_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT116), .B(new_n751_), .C1(new_n744_), .C2(new_n398_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n750_), .A3(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n605_), .A2(new_n755_), .A3(new_n579_), .A4(new_n691_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n603_), .A2(new_n579_), .A3(new_n593_), .A4(new_n604_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT54), .B1(new_n757_), .B2(new_n551_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n537_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n530_), .A2(KEYINPUT55), .A3(new_n531_), .A4(new_n536_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n765_), .A2(KEYINPUT118), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n530_), .A2(new_n536_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n765_), .A2(KEYINPUT118), .B1(new_n767_), .B2(new_n538_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n537_), .A2(KEYINPUT117), .A3(new_n761_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n764_), .A2(new_n766_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n546_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n770_), .A2(KEYINPUT119), .A3(new_n775_), .A4(new_n546_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n541_), .A2(new_n546_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .A4(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n566_), .A2(new_n574_), .A3(new_n569_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n567_), .A2(new_n568_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n562_), .A2(new_n565_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n568_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n783_), .B2(new_n574_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n547_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n516_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT121), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n517_), .B1(new_n779_), .B2(new_n786_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n791_), .A2(KEYINPUT57), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n784_), .B1(new_n771_), .B2(KEYINPUT56), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n771_), .A2(KEYINPUT56), .B1(new_n541_), .B2(new_n546_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n795_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n798_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT58), .A3(new_n796_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n799_), .A2(new_n648_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n648_), .A3(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT120), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n793_), .A2(new_n794_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n760_), .B1(new_n807_), .B2(new_n721_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n614_), .A2(new_n374_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n412_), .A2(new_n430_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813_), .B2(new_n692_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n816_));
  INV_X1    g615(.A(new_n811_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n802_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n593_), .B1(new_n818_), .B2(new_n794_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(new_n817_), .C1(new_n819_), .C2(new_n760_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n820_), .A2(KEYINPUT122), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(KEYINPUT122), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n815_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n579_), .A2(new_n343_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT123), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n814_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  NAND4_X1  g625(.A1(new_n815_), .A2(new_n821_), .A3(new_n551_), .A4(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n691_), .B2(G120gat), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n813_), .B(new_n830_), .C1(new_n829_), .C2(G120gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n813_), .B2(new_n593_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n593_), .A2(G127gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n823_), .B2(new_n834_), .ZN(G1342gat));
  AOI21_X1  g634(.A(G134gat), .B1(new_n813_), .B2(new_n517_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n648_), .A2(G134gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n823_), .B2(new_n837_), .ZN(G1343gat));
  INV_X1    g637(.A(new_n808_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(new_n412_), .A3(new_n448_), .A4(new_n809_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n579_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n324_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n691_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n325_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n840_), .A2(new_n721_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  NOR3_X1   g646(.A1(new_n840_), .A2(new_n334_), .A3(new_n649_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n334_), .B1(new_n840_), .B2(new_n516_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT124), .B(new_n334_), .C1(new_n840_), .C2(new_n516_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(G1347gat));
  NOR2_X1   g652(.A1(new_n615_), .A2(new_n373_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n631_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n412_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n692_), .B(new_n856_), .C1(new_n819_), .C2(new_n760_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n857_), .A2(new_n858_), .A3(G169gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n857_), .B2(G169gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n792_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT121), .B1(new_n791_), .B2(KEYINPUT57), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n794_), .B(new_n805_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n760_), .B1(new_n863_), .B2(new_n721_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n867_), .B(new_n856_), .C1(new_n819_), .C2(new_n760_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n692_), .A2(new_n225_), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n859_), .A2(new_n860_), .B1(new_n869_), .B2(new_n870_), .ZN(G1348gat));
  INV_X1    g670(.A(new_n869_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G176gat), .B1(new_n872_), .B2(new_n551_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n808_), .A2(new_n412_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n855_), .A2(new_n221_), .A3(new_n691_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n855_), .A2(new_n721_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G183gat), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n721_), .A2(new_n247_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n872_), .B2(new_n879_), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n866_), .A2(new_n648_), .A3(new_n868_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G190gat), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n866_), .A2(new_n868_), .A3(new_n244_), .A4(new_n517_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT126), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n882_), .A2(new_n886_), .A3(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1351gat));
  NOR3_X1   g687(.A1(new_n808_), .A2(new_n411_), .A3(new_n631_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n692_), .A3(new_n854_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n854_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n258_), .A2(KEYINPUT127), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n892_), .A2(new_n691_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n892_), .B2(new_n691_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1353gat));
  NAND3_X1  g695(.A1(new_n889_), .A2(new_n593_), .A3(new_n854_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT63), .B(G211gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n897_), .B2(new_n900_), .ZN(G1354gat));
  INV_X1    g700(.A(G218gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n892_), .A2(new_n902_), .A3(new_n649_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n892_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n517_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(new_n905_), .ZN(G1355gat));
endmodule


