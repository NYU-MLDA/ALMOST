//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  XNOR2_X1  g000(.A(KEYINPUT18), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT93), .ZN(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(G204gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(G197gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT21), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n211_), .B(KEYINPUT92), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(G197gat), .B2(new_n212_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n209_), .B(new_n214_), .C1(new_n216_), .C2(KEYINPUT21), .ZN(new_n217_));
  INV_X1    g016(.A(new_n209_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n216_), .A3(KEYINPUT21), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT24), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  MUX2_X1   g024(.A(new_n224_), .B(KEYINPUT24), .S(new_n225_), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT23), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n226_), .A2(new_n230_), .A3(new_n234_), .A4(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n228_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(G183gat), .B2(G190gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n222_), .A2(new_n223_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n242_), .B2(new_n223_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT95), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n221_), .A2(new_n238_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G226gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT19), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n231_), .A2(KEYINPUT81), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT25), .Z(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n252_), .A2(new_n232_), .A3(KEYINPUT26), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n252_), .B2(new_n235_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n239_), .B(new_n226_), .C1(new_n251_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n230_), .A2(new_n234_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n243_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n220_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n246_), .A2(KEYINPUT20), .A3(new_n249_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n245_), .A2(new_n238_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n220_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n220_), .A2(new_n259_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n249_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n207_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n266_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n248_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n207_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n261_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G1gat), .B(G29gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n280_), .A2(new_n281_), .B1(KEYINPUT87), .B2(KEYINPUT3), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  OAI22_X1  g085(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n282_), .A2(new_n285_), .A3(new_n286_), .A4(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n289_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n292_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT88), .A3(new_n290_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n288_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT89), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n295_), .A2(new_n293_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n288_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n303_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n290_), .A2(KEYINPUT1), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT86), .B1(new_n308_), .B2(new_n292_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n291_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n294_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n283_), .B(KEYINPUT85), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n280_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n301_), .A2(new_n306_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT96), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n314_), .A2(new_n280_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n320_), .A2(new_n315_), .B1(new_n300_), .B2(new_n297_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n304_), .A2(new_n322_), .A3(new_n305_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT84), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT96), .B1(new_n321_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n319_), .B1(new_n326_), .B2(new_n317_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n325_), .B1(new_n301_), .B2(new_n316_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(KEYINPUT4), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n321_), .A2(KEYINPUT96), .A3(new_n306_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n301_), .A2(new_n316_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n325_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n318_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n317_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n338_), .B2(KEYINPUT4), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n279_), .B(new_n330_), .C1(new_n339_), .C2(new_n329_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT99), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n317_), .B1(new_n331_), .B2(new_n318_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(new_n333_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n328_), .B1(new_n345_), .B2(new_n332_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n346_), .A2(KEYINPUT99), .A3(new_n279_), .A4(new_n330_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n273_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n345_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n338_), .A2(new_n328_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n278_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT98), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT33), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n332_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n329_), .B(new_n355_), .C1(new_n327_), .C2(new_n343_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n279_), .B1(new_n356_), .B2(new_n350_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n357_), .A2(KEYINPUT98), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n348_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT100), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n279_), .A3(new_n350_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n352_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n221_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT20), .A3(new_n260_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n248_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n248_), .B2(new_n269_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n270_), .A2(new_n261_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n364_), .B(new_n370_), .C1(new_n371_), .C2(new_n369_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n348_), .B(KEYINPUT100), .C1(new_n354_), .C2(new_n359_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n362_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n325_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(new_n259_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G15gat), .B(G43gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT31), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n376_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n379_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n334_), .A2(KEYINPUT29), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT91), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n220_), .B1(new_n385_), .B2(KEYINPUT91), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n321_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n221_), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n388_), .A2(new_n389_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT28), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n334_), .A2(KEYINPUT29), .ZN(new_n396_));
  XOR2_X1   g195(.A(G22gat), .B(G50gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT90), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n395_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(new_n401_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n374_), .A2(new_n384_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n364_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n207_), .B(KEYINPUT101), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n368_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT27), .A3(new_n272_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n273_), .A2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n402_), .A2(new_n383_), .A3(new_n403_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n383_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n406_), .B(new_n412_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n405_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G190gat), .B(G218gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G134gat), .ZN(new_n418_));
  INV_X1    g217(.A(G162gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT36), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(KEYINPUT66), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n425_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(KEYINPUT66), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n424_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT10), .B(G99gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT65), .B(G85gat), .ZN(new_n436_));
  INV_X1    g235(.A(G92gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n439_));
  INV_X1    g238(.A(KEYINPUT9), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n438_), .A2(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  OAI221_X1 g242(.A(new_n434_), .B1(G106gat), .B2(new_n435_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n445_));
  NOR2_X1   g244(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n448_), .B(new_n449_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n430_), .A2(new_n433_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n445_), .B1(new_n451_), .B2(KEYINPUT68), .ZN(new_n452_));
  INV_X1    g251(.A(new_n443_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n441_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n447_), .A2(new_n450_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n431_), .A2(new_n432_), .A3(new_n424_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n424_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n455_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n452_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT69), .B1(new_n457_), .B2(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n430_), .A2(new_n464_), .A3(new_n433_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n465_), .A3(new_n456_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n445_), .B1(new_n466_), .B2(new_n455_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n444_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469_));
  OR2_X1    g268(.A1(G29gat), .A2(G36gat), .ZN(new_n470_));
  INV_X1    g269(.A(G43gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G29gat), .A2(G36gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G50gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G43gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(G50gat), .B1(new_n479_), .B2(new_n473_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n469_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n475_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(G50gat), .A3(new_n473_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT15), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n468_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n477_), .A2(new_n480_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(new_n444_), .C1(new_n462_), .C2(new_n467_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT72), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT34), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n491_), .A2(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n488_), .B2(KEYINPUT73), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n494_), .A2(new_n496_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n423_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT75), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n488_), .A2(new_n493_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n488_), .A2(KEYINPUT73), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n501_), .B(new_n486_), .C1(new_n502_), .C2(new_n495_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n494_), .A2(new_n496_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n503_), .A2(new_n421_), .A3(new_n504_), .A4(new_n420_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT75), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n506_), .B(new_n423_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT102), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n416_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n510_), .B(KEYINPUT103), .Z(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n466_), .A2(new_n455_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n454_), .B1(new_n451_), .B2(KEYINPUT68), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT8), .B1(new_n459_), .B2(new_n460_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n520_), .A2(KEYINPUT8), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n442_), .A2(new_n443_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n434_), .B1(G106gat), .B2(new_n435_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT71), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n444_), .B(new_n518_), .C1(new_n462_), .C2(new_n467_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT70), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n520_), .A2(KEYINPUT8), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n521_), .A2(new_n522_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n518_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n468_), .A2(new_n536_), .A3(new_n519_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n528_), .A2(new_n530_), .A3(new_n535_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n527_), .A2(KEYINPUT12), .A3(new_n529_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT12), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n468_), .A2(new_n543_), .A3(new_n519_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n539_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G120gat), .B(G148gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n212_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n223_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n541_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT13), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT13), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n551_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n222_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n210_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT78), .ZN(new_n563_));
  INV_X1    g362(.A(G1gat), .ZN(new_n564_));
  INV_X1    g363(.A(G15gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT76), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G15gat), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n566_), .A2(new_n568_), .A3(G22gat), .ZN(new_n569_));
  AOI21_X1  g368(.A(G22gat), .B1(new_n566_), .B2(new_n568_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT77), .B(G8gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT14), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n564_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(G22gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n567_), .A2(G15gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n565_), .A2(KEYINPUT76), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n575_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT14), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n568_), .A3(G22gat), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n564_), .A4(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n574_), .A2(new_n582_), .A3(G8gat), .ZN(new_n583_));
  INV_X1    g382(.A(G8gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G1gat), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n586_), .B2(new_n581_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n487_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n583_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G8gat), .B1(new_n574_), .B2(new_n582_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n584_), .A3(new_n581_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n487_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n563_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n588_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n591_), .A3(new_n487_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT78), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n593_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n485_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n594_), .B(KEYINPUT79), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n596_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n599_), .A2(new_n596_), .A3(KEYINPUT80), .A4(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n562_), .B1(new_n598_), .B2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n593_), .A2(G229gat), .A3(G233gat), .A4(new_n597_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n562_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n603_), .A3(new_n604_), .A4(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n590_), .A2(new_n591_), .ZN(new_n612_));
  AND2_X1   g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n519_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT16), .B(G183gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  INV_X1    g420(.A(KEYINPUT17), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n614_), .A2(new_n615_), .A3(new_n518_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n617_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n621_), .B(new_n622_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n559_), .A2(new_n611_), .A3(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n511_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n364_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G1gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n420_), .A2(new_n421_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n497_), .A2(new_n498_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n422_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT37), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT74), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n500_), .A2(new_n640_), .A3(new_n505_), .A4(new_n507_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT74), .B(KEYINPUT37), .C1(new_n635_), .C2(new_n636_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n405_), .B2(new_n415_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(new_n630_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n564_), .A3(new_n364_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(KEYINPUT104), .A2(KEYINPUT38), .ZN(new_n648_));
  AND2_X1   g447(.A1(KEYINPUT104), .A2(KEYINPUT38), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n633_), .B(new_n650_), .C1(new_n648_), .C2(new_n647_), .ZN(G1324gat));
  INV_X1    g450(.A(new_n412_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n511_), .A2(new_n630_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(G8gat), .A3(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n646_), .A2(new_n572_), .A3(new_n652_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n656_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n653_), .A2(G8gat), .A3(new_n659_), .A4(new_n654_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n657_), .A2(KEYINPUT40), .A3(new_n658_), .A4(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1325gat));
  NAND3_X1  g464(.A1(new_n646_), .A2(new_n565_), .A3(new_n383_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n631_), .A2(new_n383_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(new_n667_), .B2(G15gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(G1326gat));
  INV_X1    g469(.A(new_n404_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n646_), .A2(new_n575_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n631_), .A2(new_n671_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G22gat), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT42), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT42), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(G1327gat));
  AOI21_X1  g476(.A(new_n509_), .B1(new_n405_), .B2(new_n415_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n559_), .A2(new_n611_), .A3(new_n628_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n364_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n416_), .A2(new_n644_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n416_), .A2(new_n684_), .A3(new_n644_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT106), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT106), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n686_), .A2(new_n679_), .A3(new_n688_), .A4(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n684_), .B1(new_n416_), .B2(new_n644_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n643_), .C1(new_n405_), .C2(new_n415_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n679_), .B(new_n688_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n689_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n406_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n681_), .B1(new_n696_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n680_), .A2(new_n698_), .A3(new_n652_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT45), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n694_), .A2(new_n689_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n694_), .A2(new_n689_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n652_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n704_), .B2(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n412_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n706_), .A2(KEYINPUT107), .A3(new_n698_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n700_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT46), .B(new_n700_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  NAND3_X1  g511(.A1(new_n680_), .A2(new_n471_), .A3(new_n383_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n384_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n471_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n680_), .B2(new_n671_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n404_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G50gat), .ZN(G1331gat));
  NAND2_X1  g518(.A1(new_n611_), .A2(new_n628_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n558_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n511_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT109), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n511_), .A2(new_n724_), .A3(new_n721_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n723_), .A2(G57gat), .A3(new_n364_), .A4(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n645_), .A2(new_n721_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n364_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT108), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1332gat));
  NOR2_X1   g529(.A1(new_n412_), .A2(G64gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT110), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n723_), .A2(new_n652_), .A3(new_n725_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G64gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G64gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1333gat));
  NOR2_X1   g537(.A1(new_n384_), .A2(G71gat), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n727_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n723_), .A2(new_n383_), .A3(new_n725_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(G71gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G71gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n727_), .A2(new_n747_), .A3(new_n671_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n723_), .A2(new_n671_), .A3(new_n725_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G78gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G78gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1335gat));
  NOR3_X1   g552(.A1(new_n558_), .A2(new_n610_), .A3(new_n628_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n678_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n364_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n686_), .A2(new_n754_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n406_), .A2(new_n436_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n755_), .B2(new_n652_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n412_), .A2(new_n437_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n757_), .B2(new_n761_), .ZN(G1337gat));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n383_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n384_), .A2(new_n435_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n763_), .A2(G99gat), .B1(new_n755_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n767_), .B(new_n768_), .Z(G1338gat));
  NAND3_X1  g568(.A1(new_n755_), .A2(new_n449_), .A3(new_n671_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n757_), .A2(new_n671_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G106gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT52), .B(new_n449_), .C1(new_n757_), .C2(new_n671_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  OAI21_X1  g576(.A(G113gat), .B1(new_n611_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n413_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n593_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n599_), .A2(new_n596_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n780_), .B(new_n562_), .C1(new_n781_), .C2(new_n600_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n609_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n552_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n542_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n545_), .B2(new_n539_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT55), .B(new_n540_), .C1(new_n542_), .C2(new_n544_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n785_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n550_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n790_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n784_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n643_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT58), .B(new_n784_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT115), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  INV_X1    g597(.A(new_n785_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n546_), .A2(KEYINPUT55), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n545_), .A2(new_n786_), .A3(new_n539_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n802_), .B2(new_n550_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n790_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT58), .A4(new_n784_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n795_), .A2(new_n797_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n783_), .B1(new_n555_), .B2(new_n551_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n610_), .A2(KEYINPUT114), .A3(new_n551_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT114), .B1(new_n610_), .B2(new_n551_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n805_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT102), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n508_), .B(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n809_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n810_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n791_), .A2(new_n792_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n610_), .A2(new_n551_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n610_), .A2(KEYINPUT114), .A3(new_n551_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n509_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n808_), .A2(new_n817_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n629_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n720_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n643_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT54), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n643_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT113), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n832_), .B(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n779_), .B1(new_n828_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n652_), .A2(new_n406_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n842_), .B(new_n840_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n843_));
  OAI221_X1 g642(.A(new_n778_), .B1(new_n777_), .B2(G113gat), .C1(new_n841_), .C2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n838_), .A2(new_n610_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(G113gat), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n844_), .A2(KEYINPUT118), .A3(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n841_), .A2(new_n843_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT120), .B1(new_n852_), .B2(new_n558_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT119), .B(G120gat), .Z(new_n854_));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n559_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n558_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n838_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1341gat));
  AOI21_X1  g660(.A(G127gat), .B1(new_n838_), .B2(new_n628_), .ZN(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n852_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n864_), .B2(new_n628_), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n838_), .B2(new_n816_), .ZN(new_n866_));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n852_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n868_), .B2(new_n644_), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n828_), .A2(new_n835_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(new_n414_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n837_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n610_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n559_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n872_), .A2(new_n629_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  OAI21_X1  g679(.A(new_n419_), .B1(new_n872_), .B2(new_n509_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n644_), .A2(G162gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT121), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n872_), .B2(new_n883_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT122), .Z(G1347gat));
  NOR2_X1   g684(.A1(new_n412_), .A2(new_n364_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n870_), .A2(new_n610_), .A3(new_n413_), .A4(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT123), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n836_), .A2(new_n889_), .A3(new_n610_), .A4(new_n886_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(G169gat), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n888_), .A2(KEYINPUT124), .A3(G169gat), .A4(new_n890_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(KEYINPUT62), .A3(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n610_), .A2(KEYINPUT125), .A3(new_n242_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  INV_X1    g696(.A(new_n242_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n611_), .B2(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n836_), .A2(new_n896_), .A3(new_n886_), .A4(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n891_), .A2(new_n892_), .A3(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n895_), .A2(new_n900_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT126), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n895_), .A2(new_n905_), .A3(new_n900_), .A4(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1348gat));
  NAND2_X1  g706(.A1(new_n836_), .A2(new_n886_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n558_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n223_), .ZN(G1349gat));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n629_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n236_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n231_), .B2(new_n911_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n908_), .B2(new_n643_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n816_), .A2(new_n235_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n908_), .B2(new_n915_), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n871_), .A2(new_n886_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n611_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n210_), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n558_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n212_), .ZN(G1353gat));
  NAND3_X1  g720(.A1(new_n871_), .A2(new_n628_), .A3(new_n886_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n923_), .ZN(G1354gat));
  NOR2_X1   g725(.A1(new_n917_), .A2(new_n509_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n644_), .A2(G218gat), .ZN(new_n928_));
  OAI22_X1  g727(.A1(new_n927_), .A2(G218gat), .B1(new_n917_), .B2(new_n928_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


