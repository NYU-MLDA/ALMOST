//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n211_), .C1(new_n212_), .C2(KEYINPUT64), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(KEYINPUT64), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT10), .B(G99gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(G106gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT65), .B1(new_n215_), .B2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n226_), .A2(new_n227_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n228_), .B(new_n229_), .C1(new_n214_), .C2(new_n213_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n210_), .A2(KEYINPUT66), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n227_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  AOI211_X1 g036(.A(KEYINPUT8), .B(new_n232_), .C1(new_n237_), .C2(new_n220_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n220_), .A2(new_n236_), .A3(new_n235_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n232_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n223_), .B(new_n230_), .C1(new_n238_), .C2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G29gat), .B(G36gat), .Z(new_n244_));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  OR2_X1    g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT75), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n246_), .B(KEYINPUT15), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n223_), .A2(new_n230_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n241_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT8), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n240_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n247_), .B(new_n248_), .C1(new_n249_), .C2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n207_), .B1(new_n258_), .B2(KEYINPUT74), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n248_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n249_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n256_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n250_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n260_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266_));
  INV_X1    g065(.A(new_n207_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT34), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n259_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n259_), .B2(new_n268_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n206_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n259_), .A2(new_n268_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n271_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n205_), .B(KEYINPUT36), .Z(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(G43gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(G15gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n283_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT25), .B(G183gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n291_));
  OR2_X1    g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT24), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT23), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(KEYINPUT24), .B2(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n294_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(KEYINPUT81), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G169gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(G176gat), .B1(new_n302_), .B2(KEYINPUT82), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT22), .B(G169gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(KEYINPUT82), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT83), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n303_), .B(new_n307_), .C1(KEYINPUT82), .C2(new_n304_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n293_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n296_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n295_), .A2(new_n300_), .B1(new_n309_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n309_), .A2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n299_), .A2(KEYINPUT81), .ZN(new_n320_));
  INV_X1    g119(.A(new_n298_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n295_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n319_), .A2(new_n322_), .A3(new_n317_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n318_), .A2(new_n323_), .A3(KEYINPUT85), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT85), .B1(new_n318_), .B2(new_n323_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n287_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n325_), .A2(new_n287_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G134gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT31), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OR3_X1    g131(.A1(new_n326_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n332_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G141gat), .B(G148gat), .Z(new_n337_));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT86), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT1), .ZN(new_n340_));
  OR2_X1    g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n340_), .B(new_n341_), .C1(KEYINPUT1), .C2(new_n338_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n339_), .B1(new_n338_), .B2(KEYINPUT1), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n337_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  INV_X1    g144(.A(G141gat), .ZN(new_n346_));
  INV_X1    g145(.A(G148gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n344_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT87), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n344_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n358_), .A3(new_n330_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n355_), .A2(new_n330_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n360_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n356_), .A2(new_n364_), .A3(new_n358_), .A4(new_n330_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n362_), .B1(new_n363_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT95), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G85gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT94), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n363_), .A2(new_n367_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n362_), .A2(new_n373_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n365_), .A2(new_n366_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n360_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n383_), .A3(KEYINPUT94), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n368_), .A2(new_n374_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n379_), .A2(new_n384_), .B1(new_n385_), .B2(KEYINPUT95), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387_));
  OR2_X1    g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT21), .A3(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G211gat), .B(G218gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT89), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT21), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT88), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n397_), .A3(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n391_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n392_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  AOI211_X1 g201(.A(KEYINPUT89), .B(new_n400_), .C1(new_n396_), .C2(new_n398_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n356_), .A2(new_n358_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n387_), .B(new_n404_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(new_n401_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n392_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n355_), .A2(KEYINPUT29), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n413_));
  INV_X1    g212(.A(new_n398_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n397_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n401_), .B(new_n413_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n387_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n400_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n420_), .B2(new_n392_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n344_), .B2(new_n354_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n408_), .B(new_n418_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n407_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n344_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n357_), .B1(new_n344_), .B2(new_n354_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT28), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n405_), .A2(new_n432_), .A3(new_n406_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G22gat), .B(G50gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n431_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n426_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n407_), .C1(new_n419_), .C2(new_n424_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n427_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n427_), .B2(new_n440_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n375_), .B(new_n386_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n297_), .B1(G183gat), .B2(G190gat), .ZN(new_n445_));
  INV_X1    g244(.A(G176gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n310_), .B1(new_n304_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n299_), .B2(new_n298_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n444_), .B1(new_n404_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT19), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n421_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n316_), .B2(new_n421_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n299_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n321_), .A2(new_n456_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n421_), .A2(KEYINPUT91), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT91), .B1(new_n421_), .B2(new_n457_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n455_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n454_), .B1(new_n460_), .B2(new_n452_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G8gat), .B(G36gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT18), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n452_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n319_), .A2(new_n322_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n444_), .B1(new_n469_), .B2(new_n404_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n457_), .A2(KEYINPUT93), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n449_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n473_), .A3(new_n421_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n468_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n411_), .A2(new_n416_), .A3(new_n449_), .ZN(new_n476_));
  AND4_X1   g275(.A1(KEYINPUT20), .A2(new_n453_), .A3(new_n468_), .A4(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n467_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT96), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT96), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n480_), .B(new_n467_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n466_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT27), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT27), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n467_), .B(new_n454_), .C1(new_n460_), .C2(new_n452_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n466_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n443_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n442_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n427_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n379_), .A2(new_n384_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n359_), .A2(new_n360_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n382_), .A2(new_n381_), .B1(new_n492_), .B2(new_n361_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT95), .B1(new_n493_), .B2(new_n373_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n375_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n465_), .A2(KEYINPUT32), .ZN(new_n496_));
  INV_X1    g295(.A(new_n474_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n452_), .B1(new_n497_), .B2(new_n455_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n450_), .A2(new_n468_), .A3(new_n453_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n496_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(new_n461_), .B2(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n380_), .A2(new_n383_), .A3(KEYINPUT33), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT33), .B1(new_n380_), .B2(new_n383_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n382_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n492_), .A2(new_n366_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(new_n374_), .ZN(new_n509_));
  AOI211_X1 g308(.A(KEYINPUT92), .B(new_n373_), .C1(new_n492_), .C2(new_n366_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n506_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n466_), .A3(new_n511_), .A4(new_n485_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n490_), .B1(new_n502_), .B2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT97), .B(new_n336_), .C1(new_n487_), .C2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n336_), .A2(new_n490_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n495_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n483_), .A2(new_n486_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n502_), .A2(new_n512_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n441_), .A2(new_n442_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n461_), .A2(new_n465_), .B1(new_n478_), .B2(KEYINPUT96), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n484_), .B1(new_n523_), .B2(new_n481_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n486_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n516_), .B(new_n490_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT97), .B1(new_n527_), .B2(new_n336_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT99), .B(new_n281_), .C1(new_n519_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531_));
  INV_X1    g330(.A(new_n443_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n517_), .A2(new_n532_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n533_), .B2(new_n335_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n518_), .A3(new_n514_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT99), .B1(new_n535_), .B2(new_n281_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n538_));
  INV_X1    g337(.A(G57gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(G64gat), .ZN(new_n540_));
  INV_X1    g339(.A(G64gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(G57gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n538_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(G57gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(G64gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT67), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G71gat), .B(G78gat), .Z(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n547_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT11), .ZN(new_n553_));
  AOI211_X1 g352(.A(KEYINPUT68), .B(new_n544_), .C1(new_n543_), .C2(new_n547_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT67), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT67), .B1(new_n545_), .B2(new_n546_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT11), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT68), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n551_), .A3(KEYINPUT11), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n548_), .A4(new_n549_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n243_), .A2(new_n555_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n243_), .B1(new_n561_), .B2(new_n555_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n555_), .A2(new_n561_), .A3(KEYINPUT12), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n264_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n555_), .A2(new_n561_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n243_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(new_n562_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G176gat), .B(G204gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT71), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT72), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n574_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT13), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G15gat), .B(G22gat), .ZN(new_n589_));
  INV_X1    g388(.A(G8gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G1gat), .B(G8gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n570_), .B(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n599_));
  XOR2_X1   g398(.A(G127gat), .B(G155gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n598_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n261_), .A2(new_n594_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n246_), .A2(new_n594_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n246_), .B(new_n594_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n611_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n609_), .A2(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT79), .ZN(new_n617_));
  XOR2_X1   g416(.A(G169gat), .B(G197gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n615_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n588_), .A2(new_n608_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n537_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n202_), .B1(new_n623_), .B2(new_n495_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n519_), .A2(new_n528_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n588_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n608_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n276_), .A2(new_n280_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n279_), .B(KEYINPUT76), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n278_), .A2(new_n273_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n628_), .B1(new_n276_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT77), .B1(new_n629_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n276_), .A2(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT37), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT77), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n276_), .A2(new_n280_), .A3(new_n628_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n626_), .A2(new_n627_), .A3(new_n634_), .A4(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n620_), .B(KEYINPUT80), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n625_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n495_), .A2(KEYINPUT98), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n495_), .A2(KEYINPUT98), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(new_n202_), .A3(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT38), .Z(new_n649_));
  NOR2_X1   g448(.A1(new_n624_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT100), .ZN(G1324gat));
  INV_X1    g450(.A(new_n517_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n643_), .A2(new_n590_), .A3(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n652_), .B(new_n622_), .C1(new_n530_), .C2(new_n536_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G8gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT101), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(new_n658_), .A3(G8gat), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n656_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n653_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n653_), .B(new_n663_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  NAND3_X1  g466(.A1(new_n643_), .A2(new_n285_), .A3(new_n335_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n537_), .A2(new_n335_), .A3(new_n622_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n669_), .B2(G15gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n643_), .A2(new_n674_), .A3(new_n490_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n623_), .A2(new_n490_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G22gat), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT42), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT42), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1327gat));
  NOR2_X1   g479(.A1(new_n625_), .A2(new_n642_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n588_), .A2(new_n281_), .A3(new_n627_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n495_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n634_), .A2(new_n639_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n519_), .B2(new_n528_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n535_), .A2(KEYINPUT43), .A3(new_n686_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n588_), .A2(new_n621_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n689_), .A2(new_n690_), .A3(new_n608_), .A4(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n696_), .A3(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n689_), .A2(new_n608_), .A3(new_n690_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(KEYINPUT106), .A3(KEYINPUT44), .A4(new_n691_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n627_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n701_), .A2(KEYINPUT44), .A3(new_n691_), .A4(new_n690_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n698_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n647_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n685_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n702_), .A2(new_n703_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n702_), .A2(new_n703_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n652_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n697_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n696_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G36gat), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n683_), .A2(G36gat), .A3(new_n517_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n709_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n517_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n698_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n709_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n723_), .A2(new_n718_), .A3(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n720_), .A2(new_n725_), .ZN(G1329gat));
  NAND4_X1  g525(.A1(new_n698_), .A2(new_n705_), .A3(G43gat), .A4(new_n335_), .ZN(new_n727_));
  INV_X1    g526(.A(G43gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n683_), .B2(new_n336_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n727_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n684_), .B2(new_n490_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n490_), .A2(G50gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n706_), .B2(new_n735_), .ZN(G1331gat));
  NOR3_X1   g535(.A1(new_n626_), .A2(new_n608_), .A3(new_n641_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n537_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n516_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n535_), .A2(new_n621_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n626_), .B1(new_n741_), .B2(KEYINPUT109), .ZN(new_n742_));
  OR3_X1    g541(.A1(new_n625_), .A2(KEYINPUT109), .A3(new_n620_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n686_), .A2(new_n608_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n539_), .A3(new_n647_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n740_), .A2(new_n747_), .ZN(G1332gat));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n541_), .A3(new_n652_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G64gat), .B1(new_n739_), .B2(new_n517_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT48), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT48), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n754_), .A3(new_n335_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G71gat), .B1(new_n739_), .B2(new_n336_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT49), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT49), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(G1334gat));
  INV_X1    g558(.A(G78gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n746_), .A2(new_n760_), .A3(new_n490_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n738_), .A2(new_n490_), .ZN(new_n762_));
  XOR2_X1   g561(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(G78gat), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n626_), .A2(new_n620_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n699_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT111), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n699_), .A2(new_n770_), .A3(new_n767_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n516_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n627_), .A2(new_n281_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n744_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n208_), .A3(new_n647_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1336gat));
  OAI21_X1  g576(.A(G92gat), .B1(new_n772_), .B2(new_n517_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n209_), .A3(new_n652_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1337gat));
  NOR2_X1   g579(.A1(new_n336_), .A2(new_n221_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n744_), .A2(new_n774_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT51), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n336_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(new_n234_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n783_), .A2(KEYINPUT51), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n699_), .A2(new_n490_), .A3(new_n767_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT114), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n792_), .A2(KEYINPUT52), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(KEYINPUT114), .A3(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n521_), .A2(G106gat), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n742_), .A2(new_n743_), .A3(new_n774_), .A4(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n797_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT53), .B1(new_n795_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n792_), .A2(KEYINPUT52), .A3(new_n794_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n797_), .A4(new_n801_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1339gat));
  NAND3_X1  g606(.A1(new_n647_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n555_), .A2(new_n561_), .A3(KEYINPUT12), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n257_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n572_), .A2(KEYINPUT12), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n562_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n566_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n565_), .A2(KEYINPUT55), .A3(new_n566_), .A4(new_n568_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n566_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n569_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n581_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n809_), .B(KEYINPUT56), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n582_), .A2(new_n620_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n818_), .A2(new_n822_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT116), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n581_), .A3(new_n823_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n809_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT118), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n809_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n826_), .A4(new_n827_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n609_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n619_), .B1(new_n613_), .B2(new_n611_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n615_), .A2(new_n619_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n584_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n833_), .A2(new_n838_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n281_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n831_), .A2(KEYINPUT56), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n830_), .A2(new_n835_), .A3(new_n581_), .A4(new_n823_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n582_), .A2(new_n841_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n848_), .A2(KEYINPUT58), .A3(new_n849_), .A4(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n686_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n847_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n843_), .B2(new_n281_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n608_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n640_), .B2(new_n641_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n745_), .A2(new_n861_), .A3(new_n626_), .A4(new_n642_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n808_), .B1(new_n859_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n620_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT119), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n865_), .A2(new_n869_), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT120), .B1(new_n864_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n860_), .A2(new_n862_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n843_), .A2(new_n281_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n845_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n843_), .A2(new_n846_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n879_), .B2(new_n608_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n874_), .B(KEYINPUT59), .C1(new_n880_), .C2(new_n808_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n873_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n808_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n627_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n872_), .B(new_n883_), .C1(new_n884_), .C2(new_n875_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n859_), .A2(new_n863_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(KEYINPUT121), .A3(new_n872_), .A4(new_n883_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n882_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n642_), .A2(new_n866_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n871_), .B1(new_n891_), .B2(new_n892_), .ZN(G1340gat));
  NAND3_X1  g692(.A1(new_n882_), .A2(new_n588_), .A3(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G120gat), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n864_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n896_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1341gat));
  NAND3_X1  g698(.A1(new_n882_), .A2(new_n627_), .A3(new_n890_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G127gat), .ZN(new_n901_));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n864_), .A2(new_n902_), .A3(new_n627_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1342gat));
  AOI21_X1  g703(.A(G134gat), .B1(new_n864_), .B2(new_n844_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n686_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT122), .B(G134gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n891_), .B2(new_n908_), .ZN(G1343gat));
  NOR3_X1   g708(.A1(new_n652_), .A2(new_n335_), .A3(new_n521_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n888_), .A2(new_n647_), .A3(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n621_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n346_), .ZN(G1344gat));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n626_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT123), .B(G148gat), .Z(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1345gat));
  NOR2_X1   g715(.A1(new_n911_), .A2(new_n608_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT61), .B(G155gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n911_), .B2(new_n906_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n281_), .A2(G162gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n911_), .B2(new_n921_), .ZN(G1347gat));
  NOR3_X1   g721(.A1(new_n647_), .A2(new_n336_), .A3(new_n517_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n888_), .A2(new_n521_), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924_), .B2(new_n621_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n926_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n924_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n929_), .A2(new_n304_), .A3(new_n620_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n928_), .A3(new_n930_), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n929_), .B2(new_n588_), .ZN(new_n932_));
  OR3_X1    g731(.A1(new_n880_), .A2(KEYINPUT124), .A3(new_n490_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n880_), .B2(new_n490_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n923_), .A2(G176gat), .A3(new_n588_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n932_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  NOR3_X1   g736(.A1(new_n924_), .A2(new_n288_), .A3(new_n608_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n933_), .A2(new_n627_), .A3(new_n923_), .A4(new_n934_), .ZN(new_n939_));
  INV_X1    g738(.A(G183gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n924_), .B2(new_n906_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n844_), .A2(new_n289_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n924_), .B2(new_n943_), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n652_), .A2(new_n336_), .A3(new_n532_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n880_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n620_), .ZN(new_n947_));
  INV_X1    g746(.A(G197gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(KEYINPUT125), .B2(new_n948_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT125), .B(G197gat), .Z(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n947_), .B2(new_n950_), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n946_), .A2(new_n588_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g752(.A1(new_n946_), .A2(new_n627_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(KEYINPUT63), .B(G211gat), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957_));
  INV_X1    g756(.A(G211gat), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n954_), .A2(new_n957_), .A3(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(KEYINPUT126), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n954_), .A2(new_n961_), .A3(new_n957_), .A4(new_n958_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n956_), .B1(new_n960_), .B2(new_n962_), .ZN(G1354gat));
  AOI21_X1  g762(.A(G218gat), .B1(new_n946_), .B2(new_n844_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n686_), .A2(G218gat), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(KEYINPUT127), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n964_), .B1(new_n946_), .B2(new_n966_), .ZN(G1355gat));
endmodule


