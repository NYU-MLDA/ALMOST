//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT73), .B(G8gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n202_), .B(new_n208_), .C1(new_n205_), .C2(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(KEYINPUT15), .A3(new_n216_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n220_), .A2(new_n210_), .A3(new_n211_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT75), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n218_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n212_), .A2(new_n217_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n225_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n218_), .A2(new_n230_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT76), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G169gat), .B(G197gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n232_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  AND2_X1   g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(G92gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n240_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n239_), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n252_));
  NOR2_X1   g051(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n244_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n248_), .A2(new_n249_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT66), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(G99gat), .B2(G106gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G99gat), .A2(G106gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT6), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT10), .B(G99gat), .Z(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OR3_X1    g066(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n268_), .B(new_n269_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n240_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n244_), .A2(KEYINPUT67), .A3(new_n255_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT8), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT8), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n270_), .A2(new_n275_), .A3(new_n278_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n259_), .A2(new_n267_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT35), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n280_), .A2(new_n217_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n286_));
  AOI221_X4 g085(.A(new_n239_), .B1(new_n248_), .B2(new_n249_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT66), .B1(new_n256_), .B2(new_n257_), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT69), .B(new_n267_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n277_), .A2(new_n279_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT69), .B1(new_n259_), .B2(new_n267_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n220_), .A2(new_n221_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n286_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n285_), .A2(new_n281_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OAI221_X1 g096(.A(new_n286_), .B1(new_n281_), .B2(new_n285_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G190gat), .B(G218gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G134gat), .B(G162gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT36), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n298_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT71), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n297_), .A2(new_n298_), .A3(new_n305_), .A4(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n297_), .A2(new_n298_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n301_), .B(KEYINPUT36), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n304_), .A2(new_n306_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n259_), .A2(new_n267_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n290_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G57gat), .B(G64gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G78gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT11), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(KEYINPUT11), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n321_), .A2(KEYINPUT11), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n323_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n280_), .A2(new_n328_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G230gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n333_), .B(new_n335_), .C1(new_n331_), .C2(new_n330_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(KEYINPUT12), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT12), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n280_), .B2(new_n328_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n339_), .A2(new_n334_), .A3(new_n341_), .A4(new_n332_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G120gat), .B(G148gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT5), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G176gat), .B(G204gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n336_), .A2(new_n342_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT13), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(KEYINPUT13), .A3(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G231gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT74), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n212_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(new_n328_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G127gat), .B(G155gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT16), .ZN(new_n362_));
  XOR2_X1   g161(.A(G183gat), .B(G211gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT17), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT17), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n360_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n318_), .A2(new_n356_), .A3(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G197gat), .B(G204gat), .Z(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT21), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G197gat), .B(G204gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT21), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G211gat), .B(G218gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  OR3_X1    g176(.A1(new_n373_), .A2(new_n376_), .A3(new_n374_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT87), .ZN(new_n380_));
  INV_X1    g179(.A(G228gat), .ZN(new_n381_));
  INV_X1    g180(.A(G233gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n377_), .A2(new_n378_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n390_), .A2(KEYINPUT84), .B1(new_n391_), .B2(KEYINPUT1), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n389_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G155gat), .B(G162gat), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n392_), .B(new_n396_), .C1(KEYINPUT1), .C2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n397_), .A2(KEYINPUT1), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(KEYINPUT85), .A3(new_n396_), .A4(new_n392_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n397_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT2), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n390_), .A2(KEYINPUT3), .B1(new_n407_), .B2(new_n393_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n406_), .B(new_n408_), .C1(KEYINPUT3), .C2(new_n390_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n400_), .A2(new_n402_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT88), .B1(new_n388_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n400_), .A2(new_n402_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n403_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT29), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n385_), .B(KEYINPUT87), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n384_), .A4(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT90), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n425_));
  OAI21_X1  g224(.A(new_n385_), .B1(new_n410_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n383_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n424_), .B1(new_n421_), .B2(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n410_), .A2(new_n411_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(KEYINPUT28), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(KEYINPUT28), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G22gat), .B(G50gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n429_), .A2(new_n430_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n430_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n437_), .A2(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n428_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT79), .B(G176gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT22), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G169gat), .ZN(new_n451_));
  INV_X1    g250(.A(G169gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT22), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G183gat), .A2(G190gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT23), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G169gat), .A2(G176gat), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n454_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n462_));
  INV_X1    g261(.A(G176gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n452_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n457_), .B(KEYINPUT23), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT25), .B(G183gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT26), .B(G190gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n452_), .A3(new_n463_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n465_), .A2(new_n466_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n473_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n461_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT20), .B1(new_n476_), .B2(new_n379_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n448_), .B1(new_n450_), .B2(G169gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n453_), .B(KEYINPUT78), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n459_), .B(new_n460_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n469_), .B(KEYINPUT77), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n464_), .A2(KEYINPUT24), .A3(new_n460_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n464_), .A2(KEYINPUT24), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n466_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n419_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n447_), .B1(new_n477_), .B2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n447_), .B1(new_n476_), .B2(new_n379_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n419_), .B2(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G8gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT18), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n444_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n477_), .A2(new_n489_), .A3(new_n447_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n447_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n461_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n379_), .A3(new_n472_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n493_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n500_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n509_), .B(KEYINPUT27), .C1(new_n500_), .C2(new_n495_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n443_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G43gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT81), .B(G15gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G227gat), .A2(G233gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n488_), .B(KEYINPUT30), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n521_), .B2(KEYINPUT82), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT82), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n523_), .A3(new_n519_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G127gat), .B(G134gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G120gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT31), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT83), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(KEYINPUT31), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n527_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n525_), .A2(new_n535_), .A3(new_n526_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n410_), .A2(new_n530_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G225gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n410_), .A2(new_n530_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n545_), .A2(new_n540_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n540_), .A2(new_n546_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n542_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n544_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G1gat), .B(G29gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G85gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT0), .B(G57gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n544_), .B(new_n555_), .C1(new_n547_), .C2(new_n550_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT96), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n560_), .A3(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n512_), .A2(new_n539_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n539_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n499_), .A2(KEYINPUT32), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n495_), .A2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n504_), .A2(new_n508_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n566_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n490_), .A2(new_n567_), .A3(new_n494_), .A4(new_n565_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(new_n561_), .A3(new_n559_), .A4(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n558_), .B(KEYINPUT33), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n501_), .A2(new_n502_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n545_), .B2(new_n540_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n541_), .A2(KEYINPUT94), .A3(new_n543_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n549_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n548_), .A2(new_n542_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n578_), .B(new_n556_), .C1(new_n547_), .C2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n443_), .B1(new_n572_), .B2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n503_), .A2(new_n510_), .A3(new_n439_), .A4(new_n442_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n562_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n564_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n586_));
  AOI211_X1 g385(.A(new_n238_), .B(new_n370_), .C1(new_n563_), .C2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(new_n204_), .A3(new_n584_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n315_), .B1(new_n586_), .B2(new_n563_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n355_), .A2(new_n238_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n369_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n597_), .B2(new_n562_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n588_), .A2(new_n589_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n590_), .A2(new_n598_), .A3(new_n599_), .ZN(G1324gat));
  INV_X1    g399(.A(new_n511_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G8gat), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT39), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n587_), .A2(new_n203_), .A3(new_n511_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(G1325gat));
  INV_X1    g406(.A(G15gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n596_), .B2(new_n539_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT41), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n587_), .A2(new_n608_), .A3(new_n539_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1326gat));
  INV_X1    g411(.A(G22gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n443_), .B(KEYINPUT97), .Z(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n596_), .B2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT42), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n587_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1327gat));
  NAND2_X1  g417(.A1(new_n586_), .A2(new_n563_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n315_), .A2(new_n594_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT99), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n592_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT100), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n619_), .A2(new_n624_), .A3(new_n592_), .A4(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OR3_X1    g425(.A1(new_n626_), .A2(G29gat), .A3(new_n562_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n593_), .A2(new_n369_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n619_), .B2(new_n317_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT43), .B(new_n318_), .C1(new_n586_), .C2(new_n563_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n628_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT44), .B(new_n628_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n584_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G29gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n636_), .B2(new_n584_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n627_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  NOR2_X1   g440(.A1(new_n601_), .A2(G36gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n623_), .A2(new_n625_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT101), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n623_), .A2(new_n645_), .A3(new_n625_), .A4(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n634_), .A2(new_n511_), .A3(new_n635_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(KEYINPUT45), .A3(new_n646_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n648_), .A2(new_n647_), .B1(new_n650_), .B2(G36gat), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n659_), .A2(new_n654_), .A3(new_n655_), .A4(new_n652_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1329gat));
  NOR2_X1   g460(.A1(new_n564_), .A2(new_n514_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n634_), .A2(new_n635_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT103), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n634_), .A2(new_n665_), .A3(new_n635_), .A4(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n514_), .B1(new_n626_), .B2(new_n564_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT104), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n667_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1330gat));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n636_), .A2(new_n443_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G50gat), .ZN(new_n676_));
  INV_X1    g475(.A(G50gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT106), .B(new_n677_), .C1(new_n636_), .C2(new_n443_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n614_), .A2(new_n677_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n676_), .A2(new_n678_), .B1(new_n626_), .B2(new_n679_), .ZN(G1331gat));
  NAND2_X1  g479(.A1(new_n355_), .A2(new_n238_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n594_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n591_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n562_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n317_), .A2(new_n594_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n681_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n619_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n584_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n683_), .B2(new_n511_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(new_n692_), .A3(new_n511_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n697_), .A3(new_n539_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G71gat), .B1(new_n684_), .B2(new_n564_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT107), .Z(G1334gat));
  INV_X1    g502(.A(G78gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n683_), .B2(new_n614_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT50), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n688_), .A2(new_n704_), .A3(new_n614_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1335gat));
  OR2_X1    g507(.A1(new_n630_), .A2(new_n631_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n594_), .A3(new_n687_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n562_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n619_), .A2(new_n621_), .A3(new_n687_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n242_), .A3(new_n584_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1336gat));
  OAI21_X1  g513(.A(G92gat), .B1(new_n710_), .B2(new_n601_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n243_), .A3(new_n511_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1337gat));
  NAND3_X1  g516(.A1(new_n712_), .A2(new_n266_), .A3(new_n539_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n709_), .A2(new_n594_), .A3(new_n539_), .A4(new_n687_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G99gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G99gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g523(.A1(new_n712_), .A2(new_n265_), .A3(new_n443_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n709_), .A2(new_n594_), .A3(new_n443_), .A4(new_n687_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G106gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G106gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g530(.A(KEYINPUT59), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n512_), .A2(new_n539_), .A3(new_n584_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n227_), .A2(new_n228_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n236_), .B1(new_n735_), .B2(new_n224_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n224_), .B1(new_n223_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n737_), .B2(new_n223_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n232_), .A2(new_n236_), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n351_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n334_), .A2(KEYINPUT111), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n339_), .A2(new_n332_), .A3(new_n341_), .A4(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n334_), .A2(new_n745_), .ZN(new_n746_));
  AND4_X1   g545(.A1(new_n339_), .A2(new_n332_), .A3(new_n341_), .A4(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n747_), .B2(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n342_), .A2(new_n745_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n342_), .A2(KEYINPUT110), .A3(new_n745_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n347_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n347_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n237_), .A2(new_n350_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n742_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n311_), .A2(KEYINPUT57), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT115), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n347_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n753_), .B2(new_n347_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n741_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n232_), .A2(new_n236_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n736_), .A2(new_n739_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n350_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT114), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n740_), .A2(new_n775_), .A3(new_n350_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n756_), .A2(new_n757_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n777_), .A2(KEYINPUT58), .B1(new_n316_), .B2(new_n314_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n776_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n758_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n762_), .A2(new_n769_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n760_), .B2(new_n315_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n369_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n370_), .B2(new_n237_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n686_), .A2(new_n356_), .A3(new_n238_), .A4(new_n787_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n732_), .B(new_n734_), .C1(new_n786_), .C2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n762_), .A2(new_n769_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n778_), .A2(new_n782_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n315_), .B1(new_n765_), .B2(new_n741_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT113), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n784_), .C1(new_n760_), .C2(new_n315_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n793_), .A2(new_n794_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n799_), .B2(new_n594_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n733_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n237_), .B(new_n792_), .C1(new_n801_), .C2(new_n732_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(G113gat), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n767_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT115), .B(new_n761_), .C1(new_n765_), .C2(new_n741_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n794_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n796_), .A2(new_n798_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n594_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n791_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n734_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n238_), .A2(G113gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n803_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n803_), .A2(new_n816_), .A3(KEYINPUT117), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1340gat));
  NAND2_X1  g620(.A1(new_n813_), .A2(KEYINPUT59), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(new_n792_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n355_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G120gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n805_), .A2(new_n814_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n827_));
  AOI21_X1  g626(.A(G120gat), .B1(new_n355_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT118), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n827_), .B2(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n825_), .B1(new_n826_), .B2(new_n832_), .ZN(G1341gat));
  NAND2_X1  g632(.A1(new_n823_), .A2(new_n369_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G127gat), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n594_), .A2(G127gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n826_), .B2(new_n836_), .ZN(G1342gat));
  XOR2_X1   g636(.A(KEYINPUT119), .B(G134gat), .Z(new_n838_));
  NOR2_X1   g637(.A1(new_n318_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n805_), .A2(new_n814_), .A3(new_n315_), .ZN(new_n840_));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n823_), .A2(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n539_), .A2(new_n583_), .A3(new_n562_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n800_), .B2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n796_), .A2(new_n798_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n369_), .B1(new_n847_), .B2(new_n783_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT120), .B(new_n844_), .C1(new_n848_), .C2(new_n791_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n237_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT121), .B(G141gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n355_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n850_), .B2(new_n369_), .ZN(new_n857_));
  AOI211_X1 g656(.A(KEYINPUT122), .B(new_n594_), .C1(new_n846_), .C2(new_n849_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n857_), .A2(new_n858_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT120), .B1(new_n812_), .B2(new_n844_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n843_), .B(new_n845_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n369_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT122), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n850_), .A2(new_n856_), .A3(new_n369_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n859_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n861_), .A2(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(new_n850_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n869_), .A2(G162gat), .A3(new_n311_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G162gat), .B1(new_n869_), .B2(new_n318_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n786_), .A2(new_n791_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n539_), .A2(new_n511_), .A3(new_n562_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n614_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n237_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT124), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n873_), .A2(new_n238_), .A3(new_n875_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n452_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT62), .B1(new_n880_), .B2(new_n452_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n879_), .B1(new_n886_), .B2(new_n887_), .ZN(G1348gat));
  AOI21_X1  g687(.A(new_n448_), .B1(new_n876_), .B2(new_n355_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n800_), .A2(new_n443_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n874_), .A2(new_n356_), .A3(new_n463_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  INV_X1    g691(.A(new_n874_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n369_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(G183gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n594_), .A2(new_n467_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n876_), .B2(new_n896_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n876_), .A2(new_n315_), .A3(new_n468_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n873_), .A2(new_n318_), .A3(new_n875_), .ZN(new_n899_));
  INV_X1    g698(.A(G190gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1351gat));
  AND3_X1   g700(.A1(new_n564_), .A2(new_n443_), .A3(new_n562_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n601_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n812_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n237_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n355_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g709(.A(new_n594_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(new_n911_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n912_), .A2(KEYINPUT126), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(KEYINPUT126), .ZN(new_n914_));
  OAI22_X1  g713(.A1(new_n913_), .A2(new_n914_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n912_), .A2(KEYINPUT126), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n912_), .A2(KEYINPUT126), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n906_), .A2(new_n921_), .A3(new_n315_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n906_), .A2(new_n317_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n921_), .ZN(G1355gat));
endmodule


