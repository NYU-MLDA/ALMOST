//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(G228gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n206_), .B(KEYINPUT86), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT87), .ZN(new_n210_));
  INV_X1    g009(.A(G211gat), .ZN(new_n211_));
  INV_X1    g010(.A(G218gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT87), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G211gat), .A2(G218gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n219_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT88), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n217_), .A2(new_n220_), .A3(KEYINPUT88), .A4(new_n221_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT89), .B1(new_n217_), .B2(new_n220_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n218_), .A2(new_n219_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n228_), .A2(new_n210_), .A3(new_n229_), .A4(new_n216_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(G141gat), .B2(G148gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G141gat), .A2(G148gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT3), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n238_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n236_), .A2(KEYINPUT82), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G141gat), .A3(G148gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n246_), .A3(new_n237_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n235_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n244_), .A2(new_n246_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n241_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n233_), .A2(new_n253_), .A3(new_n234_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT29), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n208_), .B1(new_n232_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n227_), .A2(new_n230_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n255_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(new_n248_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n208_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G78gat), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n258_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n256_), .A2(KEYINPUT29), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n207_), .B1(new_n260_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n265_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n232_), .ZN(new_n272_));
  AOI21_X1  g071(.A(G78gat), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n203_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n267_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(G78gat), .A3(new_n272_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(G106gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(KEYINPUT84), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n256_), .A2(KEYINPUT29), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G22gat), .B(G50gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n281_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n278_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n274_), .A2(new_n287_), .A3(KEYINPUT84), .A4(new_n277_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G113gat), .B(G120gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G127gat), .B(G134gat), .Z(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n296_), .A2(KEYINPUT81), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT81), .B1(new_n296_), .B2(new_n298_), .ZN(new_n300_));
  OAI22_X1  g099(.A1(new_n299_), .A2(new_n300_), .B1(new_n261_), .B2(new_n248_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT95), .B1(new_n301_), .B2(KEYINPUT4), .ZN(new_n302_));
  INV_X1    g101(.A(new_n300_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(KEYINPUT81), .A3(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT95), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT4), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n256_), .A4(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n296_), .A2(new_n298_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n262_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n301_), .A3(KEYINPUT4), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT94), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n301_), .A3(KEYINPUT94), .A4(KEYINPUT4), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n309_), .A2(new_n314_), .A3(new_n316_), .A4(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n301_), .A3(new_n315_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT96), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G85gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(G1gat), .B(G29gat), .Z(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n318_), .A2(new_n320_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n305_), .A2(KEYINPUT30), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n305_), .A2(KEYINPUT30), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G169gat), .ZN(new_n333_));
  INV_X1    g132(.A(G176gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT80), .B(G176gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT22), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n337_), .B1(new_n342_), .B2(G169gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n335_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT23), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(G183gat), .B2(G190gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n335_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n333_), .A2(new_n334_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT24), .A3(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(KEYINPUT24), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n346_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT25), .B(G183gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n353_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n344_), .A2(new_n347_), .B1(new_n352_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n332_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n330_), .A2(new_n360_), .A3(new_n331_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G15gat), .B(G43gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT31), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n366_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n329_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n335_), .A2(KEYINPUT91), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n336_), .A2(new_n339_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n335_), .A2(KEYINPUT91), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT92), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT92), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n374_), .A2(new_n375_), .A3(new_n379_), .A4(new_n376_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n347_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n352_), .A2(new_n355_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n232_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT19), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n360_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n384_), .A2(KEYINPUT20), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT99), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n360_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n232_), .A2(new_n383_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n386_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n232_), .B2(new_n383_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT99), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n390_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n387_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(KEYINPUT27), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(new_n406_), .A3(new_n403_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n403_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n412_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n410_), .A2(new_n411_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n410_), .B2(new_n416_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n292_), .B(new_n373_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n421_), .A2(KEYINPUT98), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n398_), .B2(new_n420_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT98), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n329_), .B(new_n422_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n414_), .A2(new_n415_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n328_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n311_), .A2(new_n301_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n311_), .A2(new_n301_), .A3(KEYINPUT97), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n316_), .A3(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n309_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n434_));
  OAI211_X1 g233(.A(KEYINPUT33), .B(new_n433_), .C1(new_n434_), .C2(new_n316_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n325_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n321_), .A2(new_n427_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n426_), .A2(new_n428_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n425_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n329_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT27), .B1(new_n409_), .B2(new_n413_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n415_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(KEYINPUT27), .B2(new_n442_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n439_), .A2(new_n292_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n371_), .A2(new_n372_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n419_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT102), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT9), .ZN(new_n449_));
  INV_X1    g248(.A(G85gat), .ZN(new_n450_));
  INV_X1    g249(.A(G92gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n449_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n448_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G99gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT10), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT10), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G99gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(G106gat), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT64), .B(new_n455_), .C1(new_n471_), .C2(new_n449_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n457_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n458_), .A3(new_n203_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(new_n465_), .A3(new_n466_), .A4(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n478_), .B2(new_n471_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n478_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n473_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G29gat), .A2(G36gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G29gat), .A2(G36gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(G43gat), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(G29gat), .ZN(new_n486_));
  INV_X1    g285(.A(G36gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G43gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n482_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(G50gat), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(G50gat), .B1(new_n485_), .B2(new_n490_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT34), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n498_));
  OAI22_X1  g297(.A1(new_n481_), .A2(new_n495_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n485_), .A2(new_n490_), .ZN(new_n502_));
  INV_X1    g301(.A(G50gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT15), .A3(new_n491_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n481_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n497_), .A2(new_n498_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT69), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n499_), .B2(KEYINPUT70), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G190gat), .B(G218gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G134gat), .ZN(new_n514_));
  INV_X1    g313(.A(G162gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT36), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n507_), .A2(new_n511_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT71), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n512_), .A2(new_n522_), .A3(new_n519_), .A4(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n512_), .A2(new_n519_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n516_), .B(KEYINPUT36), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT101), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(KEYINPUT101), .A3(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n446_), .A2(new_n447_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n447_), .B1(new_n446_), .B2(new_n531_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G120gat), .B(G148gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n334_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(G57gat), .A2(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G57gat), .A2(G64gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT11), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n546_), .A3(new_n541_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n480_), .A2(new_n479_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n457_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n550_), .B(new_n473_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(KEYINPUT12), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n481_), .A2(new_n557_), .A3(new_n551_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT65), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n560_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT65), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n562_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n539_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT66), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n561_), .A2(new_n563_), .A3(new_n538_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n561_), .A2(KEYINPUT65), .A3(new_n563_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n566_), .B2(new_n562_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n539_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT13), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n570_), .A2(new_n579_), .A3(new_n571_), .A4(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT67), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(KEYINPUT67), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n202_), .A2(KEYINPUT72), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(G1gat), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n588_), .A3(G8gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT14), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G15gat), .B(G22gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G1gat), .B(G8gat), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n492_), .A2(new_n493_), .A3(new_n500_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT15), .B1(new_n504_), .B2(new_n491_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n595_), .B(KEYINPUT75), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n591_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n592_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n505_), .B2(new_n501_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n604_), .B2(new_n494_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n598_), .B(new_n599_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n599_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n495_), .A2(new_n595_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n604_), .A2(new_n494_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n333_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(G197gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(G197gat), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT76), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT77), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n608_), .A2(new_n612_), .A3(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n613_), .A2(KEYINPUT77), .A3(new_n619_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT16), .B(G183gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n604_), .B(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n550_), .B(KEYINPUT73), .Z(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT74), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n630_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT17), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n635_), .A3(new_n629_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT17), .B(new_n630_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n585_), .A2(new_n625_), .A3(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n534_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n202_), .B1(new_n646_), .B2(new_n329_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n524_), .A2(new_n527_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n524_), .A2(KEYINPUT37), .A3(new_n527_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n645_), .A2(new_n446_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n586_), .A2(new_n588_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n329_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n648_), .A2(new_n649_), .A3(new_n660_), .A4(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n660_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT103), .B1(new_n663_), .B2(new_n647_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1324gat));
  NOR2_X1   g464(.A1(new_n417_), .A2(new_n418_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(new_n645_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G8gat), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n667_), .A2(KEYINPUT104), .A3(G8gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT39), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G8gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n656_), .A2(new_n673_), .A3(new_n666_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n668_), .A2(new_n669_), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n674_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n674_), .A4(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1325gat));
  INV_X1    g480(.A(G15gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n656_), .A2(new_n682_), .A3(new_n445_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n646_), .A2(new_n445_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n684_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n684_), .B2(G15gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1326gat));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n291_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT105), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n656_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n646_), .A2(new_n291_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G22gat), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT42), .B(new_n688_), .C1(new_n646_), .C2(new_n291_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(new_n446_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n583_), .A2(new_n584_), .A3(new_n698_), .A4(new_n644_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n697_), .A2(new_n531_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n700_), .B2(new_n329_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n329_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n446_), .A2(new_n703_), .A3(new_n654_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n446_), .B2(new_n654_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n706_), .C2(new_n699_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n439_), .A2(new_n292_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n440_), .A2(new_n443_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n445_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n419_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n654_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT43), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n446_), .A2(new_n703_), .A3(new_n654_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(KEYINPUT106), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n699_), .A2(KEYINPUT106), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n702_), .B1(new_n707_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n701_), .B1(new_n719_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g519(.A1(new_n700_), .A2(new_n487_), .A3(new_n666_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT45), .ZN(new_n722_));
  INV_X1    g521(.A(new_n666_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n707_), .B2(new_n718_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n487_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n722_), .B(KEYINPUT46), .C1(new_n724_), .C2(new_n487_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1329gat));
  XOR2_X1   g528(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n730_));
  AND3_X1   g529(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n716_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n445_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G43gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n700_), .A2(new_n489_), .A3(new_n445_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n730_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n445_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n707_), .B2(new_n718_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n730_), .B(new_n735_), .C1(new_n738_), .C2(new_n489_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n700_), .B2(new_n291_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n292_), .B1(new_n707_), .B2(new_n718_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g543(.A(new_n585_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n643_), .A2(new_n625_), .ZN(new_n746_));
  NOR4_X1   g545(.A1(new_n697_), .A2(new_n745_), .A3(new_n654_), .A4(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n329_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n746_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n534_), .A2(new_n585_), .A3(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n702_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(G57gat), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n750_), .B2(new_n723_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT48), .ZN(new_n754_));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n747_), .A2(new_n755_), .A3(new_n666_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1333gat));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n534_), .A2(new_n445_), .A3(new_n585_), .A4(new_n749_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(G71gat), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n759_), .B2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n758_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n763_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT49), .A3(new_n761_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n737_), .A2(G71gat), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT109), .Z(new_n768_));
  NAND2_X1  g567(.A1(new_n747_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n766_), .A3(new_n769_), .ZN(G1334gat));
  OAI21_X1  g569(.A(G78gat), .B1(new_n750_), .B2(new_n292_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT50), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n747_), .A2(new_n267_), .A3(new_n291_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1335gat));
  INV_X1    g573(.A(new_n530_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n528_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n446_), .A2(new_n776_), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n698_), .B(new_n643_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n329_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n713_), .A2(new_n714_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(new_n329_), .A3(new_n778_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n782_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g582(.A(G92gat), .B1(new_n779_), .B2(new_n666_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT110), .Z(new_n785_));
  NAND4_X1  g584(.A1(new_n781_), .A2(G92gat), .A3(new_n666_), .A4(new_n778_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  NAND2_X1  g586(.A1(new_n459_), .A2(new_n461_), .ZN(new_n788_));
  AND4_X1   g587(.A1(new_n788_), .A2(new_n778_), .A3(new_n445_), .A4(new_n777_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n781_), .A2(new_n445_), .A3(new_n778_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT111), .B1(new_n792_), .B2(G99gat), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT51), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n791_), .B(new_n797_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n779_), .A2(new_n203_), .A3(new_n291_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n781_), .A2(new_n291_), .A3(new_n778_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g605(.A(G113gat), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n698_), .A2(KEYINPUT114), .A3(new_n571_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT114), .B1(new_n698_), .B2(new_n571_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n556_), .A2(new_n565_), .A3(new_n558_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n561_), .A2(KEYINPUT55), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n561_), .A2(KEYINPUT55), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n539_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(new_n539_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n598_), .B(new_n609_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n599_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n617_), .A3(new_n616_), .A4(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(new_n623_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n811_), .A2(new_n819_), .B1(new_n577_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n808_), .B1(new_n824_), .B2(new_n776_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826_));
  INV_X1    g625(.A(new_n571_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n625_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n815_), .A2(new_n539_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n816_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n698_), .A2(new_n571_), .A3(KEYINPUT114), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n815_), .A2(new_n539_), .A3(new_n816_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n828_), .A2(new_n831_), .A3(new_n832_), .A4(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n577_), .A2(new_n823_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .A3(new_n531_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(KEYINPUT56), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n815_), .A2(new_n839_), .A3(new_n539_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n838_), .A2(new_n823_), .A3(new_n571_), .A4(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n840_), .A2(new_n571_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(KEYINPUT58), .A3(new_n823_), .A4(new_n838_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n845_), .A3(new_n654_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n825_), .A2(new_n837_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n644_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT113), .B1(new_n581_), .B2(new_n749_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n851_), .B(new_n746_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n853_), .B2(new_n655_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n575_), .B1(new_n574_), .B2(new_n539_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT66), .B(new_n538_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n579_), .B1(new_n857_), .B2(new_n571_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n580_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n749_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n851_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n581_), .A2(KEYINPUT113), .A3(new_n749_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(new_n849_), .A3(new_n655_), .A4(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n848_), .B1(new_n854_), .B2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n666_), .A2(new_n702_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n737_), .A2(new_n291_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n807_), .B1(new_n868_), .B2(new_n625_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT116), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n807_), .C1(new_n868_), .C2(new_n625_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874_));
  INV_X1    g673(.A(new_n866_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n861_), .A2(new_n655_), .A3(new_n862_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT54), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n863_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n878_), .B2(new_n848_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n879_), .B2(new_n867_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n877_), .A2(new_n863_), .B1(new_n644_), .B2(new_n847_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  INV_X1    g681(.A(new_n867_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n875_), .A4(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n874_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n868_), .A2(new_n882_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n867_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(KEYINPUT117), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n625_), .B1(new_n885_), .B2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n873_), .B1(new_n889_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g689(.A(new_n868_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n745_), .B2(KEYINPUT60), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n893_), .C1(KEYINPUT60), .C2(new_n892_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n745_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n892_), .ZN(G1341gat));
  AOI21_X1  g695(.A(G127gat), .B1(new_n891_), .B2(new_n643_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n644_), .B1(new_n885_), .B2(new_n888_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g698(.A(G134gat), .B1(new_n891_), .B2(new_n776_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n885_), .A2(new_n888_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n654_), .A2(G134gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT118), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1343gat));
  NAND3_X1  g703(.A1(new_n866_), .A2(new_n291_), .A3(new_n737_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT119), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n865_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT120), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n865_), .A2(new_n909_), .A3(new_n906_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n698_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n585_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n643_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  AOI21_X1  g717(.A(G162gat), .B1(new_n911_), .B2(new_n776_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n655_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(G162gat), .B2(new_n920_), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n881_), .A2(new_n723_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n737_), .A2(new_n291_), .A3(new_n329_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n922_), .A2(new_n698_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G169gat), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n922_), .A2(new_n923_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n930_), .A2(new_n336_), .A3(new_n698_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n924_), .A2(G169gat), .A3(new_n926_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n931_), .A3(new_n932_), .ZN(G1348gat));
  NOR2_X1   g732(.A1(new_n929_), .A2(new_n745_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n340_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(G176gat), .B2(new_n934_), .ZN(G1349gat));
  NAND4_X1  g735(.A1(new_n922_), .A2(new_n353_), .A3(new_n643_), .A4(new_n923_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n865_), .A2(new_n666_), .A3(new_n643_), .A4(new_n923_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(G183gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT122), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n929_), .B2(new_n655_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n776_), .A2(new_n354_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n929_), .B2(new_n943_), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n440_), .A2(new_n737_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT123), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n922_), .A2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n625_), .ZN(new_n948_));
  XOR2_X1   g747(.A(new_n948_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n745_), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(G204gat), .Z(G1353gat));
  AOI21_X1  g750(.A(new_n644_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT124), .Z(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  OAI22_X1  g753(.A1(new_n947_), .A2(new_n953_), .B1(KEYINPUT125), .B2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(KEYINPUT125), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n956_), .B(KEYINPUT126), .Z(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n955_), .B(new_n958_), .ZN(G1354gat));
  NOR3_X1   g758(.A1(new_n947_), .A2(new_n212_), .A3(new_n655_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n922_), .A2(new_n776_), .A3(new_n946_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n212_), .B2(new_n961_), .ZN(G1355gat));
endmodule


