//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n202_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(KEYINPUT79), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n207_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G71gat), .B(G99gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(G43gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT77), .B(G15gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(G227gat), .A2(G233gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT24), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G183gat), .A3(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n228_), .A2(new_n230_), .B1(new_n231_), .B2(new_n224_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n230_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n224_), .A2(new_n231_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT75), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n226_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT76), .B(G176gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G169gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n227_), .A2(new_n229_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n243_), .B(new_n244_), .C1(G183gat), .C2(G190gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n245_), .A3(new_n222_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT78), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n208_), .B(new_n211_), .C1(new_n218_), .C2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n211_), .A2(new_n208_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n217_), .B(new_n252_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT31), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT31), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n248_), .A2(new_n249_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n253_), .A2(new_n251_), .A3(new_n256_), .A4(new_n258_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(G155gat), .B2(G162gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(G155gat), .A3(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n263_), .A2(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n267_), .B2(new_n266_), .ZN(new_n269_));
  OR2_X1    g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n271_), .B(KEYINPUT2), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT81), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n270_), .B2(KEYINPUT3), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(KEYINPUT3), .ZN(new_n277_));
  NOR3_X1   g076(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT81), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .A4(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G155gat), .B(G162gat), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n252_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n209_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n205_), .A2(KEYINPUT86), .A3(new_n207_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n286_), .A2(new_n273_), .A3(new_n282_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G225gat), .A2(G233gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G1gat), .B(G29gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT88), .B(KEYINPUT0), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n208_), .A2(new_n211_), .B1(new_n273_), .B2(new_n282_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n289_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n284_), .A2(KEYINPUT4), .A3(new_n288_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT87), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n298_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT92), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n302_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT87), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT92), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n298_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n290_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n307_), .A2(new_n313_), .B1(new_n314_), .B2(new_n295_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n262_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n226_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n221_), .A2(new_n225_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n237_), .B1(new_n320_), .B2(KEYINPUT84), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n246_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT21), .ZN(new_n324_));
  XOR2_X1   g123(.A(G211gat), .B(G218gat), .Z(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(KEYINPUT83), .ZN(new_n326_));
  XOR2_X1   g125(.A(G197gat), .B(G204gat), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n327_), .B1(KEYINPUT21), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n317_), .B1(new_n323_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n326_), .A2(new_n331_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n239_), .A2(new_n338_), .A3(new_n329_), .A4(new_n246_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n333_), .A2(new_n334_), .A3(new_n337_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n246_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n332_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n339_), .B(KEYINPUT20), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT91), .B1(new_n344_), .B2(new_n336_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n247_), .A2(new_n332_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n336_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n345_), .A3(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G8gat), .B(G36gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT93), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT94), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n344_), .A2(new_n336_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n346_), .A2(KEYINPUT20), .A3(new_n337_), .A4(new_n347_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n356_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n351_), .A2(new_n363_), .A3(new_n357_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n359_), .A2(KEYINPUT27), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n362_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n356_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n368_), .A2(KEYINPUT27), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n283_), .A2(KEYINPUT29), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n332_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n371_), .A2(new_n332_), .A3(new_n375_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT82), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n273_), .A2(new_n282_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT28), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n377_), .A2(new_n382_), .A3(KEYINPUT82), .A4(new_n378_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G22gat), .B(G50gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(new_n387_), .A3(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n316_), .A2(new_n370_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n306_), .A2(KEYINPUT89), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT33), .B(new_n298_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n367_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n302_), .B(new_n289_), .C1(KEYINPUT4), .C2(new_n284_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n284_), .A2(new_n288_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n399_), .B(new_n295_), .C1(new_n400_), .C2(new_n289_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .A4(new_n362_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT89), .B1(new_n306_), .B2(new_n394_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n396_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n351_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n360_), .A2(new_n361_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n307_), .A2(new_n313_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n314_), .A2(new_n295_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n393_), .B1(new_n404_), .B2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n365_), .A2(new_n315_), .A3(new_n391_), .A4(new_n369_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n262_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n392_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G229gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT71), .B(G15gat), .ZN(new_n419_));
  INV_X1    g218(.A(G22gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G1gat), .ZN(new_n422_));
  INV_X1    g221(.A(G8gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT72), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT72), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G1gat), .B(G8gat), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n429_), .A2(new_n431_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G29gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT69), .ZN(new_n436_));
  XOR2_X1   g235(.A(G43gat), .B(G50gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n433_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n426_), .A2(new_n428_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n430_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n438_), .B1(new_n442_), .B2(new_n432_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n418_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT15), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n438_), .B(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n442_), .A3(new_n432_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n439_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n417_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G113gat), .B(G141gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G169gat), .B(G197gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  NAND3_X1  g251(.A1(new_n444_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n416_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT68), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G78gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT11), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n462_));
  INV_X1    g261(.A(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT9), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT64), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n479_), .A3(new_n476_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  INV_X1    g284(.A(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n482_), .B1(new_n487_), .B2(new_n481_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n471_), .B(new_n474_), .C1(new_n484_), .C2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n475_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI211_X1 g293(.A(KEYINPUT8), .B(new_n490_), .C1(new_n494_), .C2(new_n471_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497_));
  INV_X1    g296(.A(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n473_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n469_), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n491_), .B(new_n499_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n490_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n496_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n466_), .B(new_n489_), .C1(new_n495_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n468_), .A2(new_n470_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n491_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT8), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n502_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n466_), .B1(new_n512_), .B2(new_n489_), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n506_), .A2(new_n513_), .A3(KEYINPUT66), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n513_), .B2(KEYINPUT66), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n489_), .B1(new_n495_), .B2(new_n504_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n466_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT12), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(new_n506_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT67), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n513_), .B2(KEYINPUT12), .ZN(new_n524_));
  AND4_X1   g323(.A1(new_n523_), .A2(new_n519_), .A3(KEYINPUT12), .A4(new_n520_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n522_), .B(new_n515_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n518_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n518_), .B2(new_n526_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n458_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n533_), .A2(new_n458_), .A3(new_n534_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n533_), .A2(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT68), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT13), .B1(new_n541_), .B2(new_n535_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n446_), .A2(new_n519_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n547_));
  OAI221_X1 g346(.A(KEYINPUT70), .B1(KEYINPUT35), .B2(new_n546_), .C1(new_n438_), .C2(new_n519_), .ZN(new_n548_));
  OR3_X1    g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n547_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n552_), .B(KEYINPUT36), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n549_), .B2(new_n554_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT37), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n549_), .A2(new_n554_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n560_), .B(new_n555_), .C1(new_n561_), .C2(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n433_), .A2(new_n434_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT73), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n520_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n466_), .A3(new_n568_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT17), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n571_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n571_), .A2(new_n573_), .B1(KEYINPUT17), .B2(new_n578_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n543_), .A2(new_n564_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n457_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n409_), .A2(new_n410_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n422_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT95), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n556_), .A2(new_n558_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n416_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n543_), .A2(new_n456_), .A3(new_n582_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n315_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n370_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n584_), .A2(G8gat), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n593_), .A2(new_n370_), .A3(new_n594_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n600_), .B2(new_n601_), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT39), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT39), .B1(new_n602_), .B2(new_n603_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n599_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n606_), .B(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n595_), .B2(new_n415_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT41), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n584_), .A2(G15gat), .A3(new_n415_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  OAI21_X1  g412(.A(G22gat), .B1(new_n595_), .B2(new_n393_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n391_), .A2(new_n420_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT98), .Z(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n584_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT99), .ZN(G1327gat));
  INV_X1    g418(.A(new_n408_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n586_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n403_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n397_), .A2(new_n401_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n622_), .A2(new_n368_), .A3(new_n623_), .A4(new_n395_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n391_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n413_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n415_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n392_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n582_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n592_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n543_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n456_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n457_), .A2(new_n636_), .A3(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(G29gat), .B1(new_n639_), .B2(new_n586_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n262_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n641_), .B(new_n564_), .C1(new_n642_), .C2(new_n392_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT100), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n629_), .A2(new_n645_), .A3(new_n641_), .A4(new_n564_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n416_), .B2(new_n563_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n543_), .A2(new_n456_), .A3(new_n630_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n586_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n640_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  NOR2_X1   g454(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT106), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n598_), .A2(G36gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n635_), .A2(new_n637_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT104), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n635_), .A2(new_n637_), .A3(new_n658_), .A4(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n650_), .A2(new_n652_), .A3(new_n598_), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n657_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n648_), .A2(new_n649_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n651_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n649_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n370_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n665_), .B1(new_n676_), .B2(G36gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n670_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n657_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n671_), .A2(new_n680_), .ZN(G1329gat));
  NAND3_X1  g480(.A1(new_n653_), .A2(G43gat), .A3(new_n262_), .ZN(new_n682_));
  INV_X1    g481(.A(G43gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n638_), .B2(new_n415_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n639_), .B2(new_n391_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n391_), .A2(G50gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n653_), .B2(new_n688_), .ZN(G1331gat));
  INV_X1    g488(.A(G57gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n543_), .A2(new_n456_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n629_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n582_), .B1(new_n562_), .B2(new_n559_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n690_), .B1(new_n696_), .B2(new_n315_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT107), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n593_), .A2(new_n630_), .A3(new_n692_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(new_n690_), .A3(new_n315_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n699_), .B2(new_n598_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n598_), .A2(G64gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n696_), .B2(new_n704_), .ZN(G1333gat));
  OAI21_X1  g504(.A(G71gat), .B1(new_n699_), .B2(new_n415_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT49), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n415_), .A2(G71gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n696_), .B2(new_n708_), .ZN(G1334gat));
  OR3_X1    g508(.A1(new_n696_), .A2(G78gat), .A3(new_n393_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n699_), .A2(new_n393_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G78gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT108), .Z(G1335gat));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n691_), .A2(new_n630_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n648_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n648_), .B2(new_n718_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(new_n586_), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n630_), .A2(new_n631_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n694_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n586_), .A2(new_n485_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n724_), .A2(new_n485_), .B1(new_n726_), .B2(new_n727_), .ZN(G1336gat));
  NAND2_X1  g527(.A1(new_n370_), .A2(G92gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n723_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n486_), .B1(new_n726_), .B2(new_n598_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1337gat));
  NAND2_X1  g532(.A1(new_n262_), .A2(new_n472_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT112), .B1(new_n726_), .B2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n262_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G99gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n737_), .B(new_n739_), .ZN(G1338gat));
  AND4_X1   g539(.A1(new_n473_), .A2(new_n694_), .A3(new_n391_), .A4(new_n725_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n648_), .A2(new_n391_), .A3(new_n718_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G106gat), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n695_), .B(new_n456_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n417_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n447_), .A2(new_n448_), .A3(new_n418_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n452_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n453_), .A2(new_n758_), .A3(new_n532_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n526_), .A2(KEYINPUT115), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT55), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n526_), .A2(KEYINPUT115), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n522_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n516_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT116), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n767_), .A3(new_n516_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n761_), .A2(new_n763_), .A3(new_n766_), .A4(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n530_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n530_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n759_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT118), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n563_), .B1(new_n773_), .B2(KEYINPUT58), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(KEYINPUT118), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n532_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n769_), .A2(new_n530_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n530_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n453_), .A2(new_n758_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n541_), .A2(new_n783_), .A3(new_n535_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT57), .B(new_n631_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n774_), .A2(new_n776_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n631_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT117), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n631_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n455_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n533_), .B1(new_n794_), .B2(new_n453_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n541_), .A2(new_n783_), .A3(new_n535_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n592_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n793_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n754_), .B1(new_n800_), .B2(new_n582_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n370_), .A2(new_n391_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n586_), .A3(new_n262_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n751_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n759_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT58), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n564_), .A3(new_n776_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n785_), .A2(new_n786_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n799_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n582_), .B1(new_n805_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n754_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n803_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n804_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n633_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n810_), .A2(new_n811_), .A3(new_n799_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n630_), .B1(new_n822_), .B2(new_n793_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT59), .B(new_n816_), .C1(new_n823_), .C2(new_n754_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n456_), .A2(KEYINPUT121), .ZN(new_n826_));
  MUX2_X1   g625(.A(KEYINPUT121), .B(new_n826_), .S(G113gat), .Z(new_n827_));
  AOI21_X1  g626(.A(new_n819_), .B1(new_n825_), .B2(new_n827_), .ZN(G1340gat));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n543_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G120gat), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n539_), .A2(new_n542_), .A3(KEYINPUT60), .ZN(new_n831_));
  MUX2_X1   g630(.A(new_n831_), .B(KEYINPUT60), .S(G120gat), .Z(new_n832_));
  NAND2_X1  g631(.A1(new_n818_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(G1341gat));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n804_), .A2(new_n817_), .A3(new_n835_), .A4(new_n630_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n582_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n835_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT122), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n836_), .B(new_n840_), .C1(new_n837_), .C2(new_n835_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1342gat));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n818_), .A2(new_n843_), .A3(new_n592_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n563_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n843_), .B2(new_n845_), .ZN(G1343gat));
  NAND4_X1  g645(.A1(new_n598_), .A2(new_n586_), .A3(new_n391_), .A4(new_n415_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT123), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n815_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n633_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n543_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g653(.A1(new_n849_), .A2(KEYINPUT124), .A3(new_n582_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT124), .B1(new_n849_), .B2(new_n582_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1346gat));
  OR3_X1    g659(.A1(new_n849_), .A2(G162gat), .A3(new_n631_), .ZN(new_n861_));
  OAI21_X1  g660(.A(G162gat), .B1(new_n849_), .B2(new_n563_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1347gat));
  NOR3_X1   g662(.A1(new_n598_), .A2(new_n316_), .A3(new_n391_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n815_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n633_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G169gat), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n241_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n869_), .B(new_n870_), .C1(new_n871_), .C2(new_n866_), .ZN(G1348gat));
  NAND3_X1  g671(.A1(new_n815_), .A2(new_n543_), .A3(new_n864_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n873_), .A2(G176gat), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n875_));
  INV_X1    g674(.A(new_n240_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n865_), .A2(new_n630_), .ZN(new_n882_));
  MUX2_X1   g681(.A(new_n219_), .B(G183gat), .S(new_n882_), .Z(G1350gat));
  NAND3_X1  g682(.A1(new_n865_), .A2(new_n220_), .A3(new_n592_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n865_), .A2(new_n564_), .ZN(new_n885_));
  INV_X1    g684(.A(G190gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1351gat));
  NAND2_X1  g686(.A1(new_n315_), .A2(new_n391_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n598_), .A2(new_n888_), .A3(new_n262_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT126), .B1(new_n815_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891_));
  INV_X1    g690(.A(new_n889_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n891_), .B(new_n892_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n893_));
  OAI211_X1 g692(.A(G197gat), .B(new_n633_), .C1(new_n890_), .C2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT127), .ZN(new_n895_));
  INV_X1    g694(.A(G197gat), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n890_), .A2(new_n893_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n456_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n891_), .B1(new_n801_), .B2(new_n892_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n815_), .A2(KEYINPUT126), .A3(new_n889_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(G197gat), .A4(new_n633_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n895_), .A2(new_n898_), .A3(new_n903_), .ZN(G1352gat));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n543_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  AND4_X1   g707(.A1(new_n630_), .A2(new_n901_), .A3(new_n907_), .A4(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n901_), .B2(new_n630_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1354gat));
  OR3_X1    g710(.A1(new_n897_), .A2(G218gat), .A3(new_n631_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G218gat), .B1(new_n897_), .B2(new_n563_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1355gat));
endmodule


