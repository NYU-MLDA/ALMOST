//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_c1355" written by ABC on Sun Mar 26 01:26:03 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n517_, new_n518_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n551_, new_n552_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n645_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n673_, new_n674_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n138_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n139_));
  NAND2_X1  g002(.A1(new_n138_), .A2(new_n139_), .ZN(new_n140_));
  XOR2_X1   g003(.A(G113gat), .B(G120gat), .Z(new_n141_));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n142_));
  NAND2_X1  g005(.A1(new_n141_), .A2(new_n142_), .ZN(new_n143_));
  NAND2_X1  g006(.A1(new_n140_), .A2(new_n143_), .ZN(new_n144_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n145_));
  XNOR2_X1  g008(.A(new_n145_), .B(KEYINPUT3), .ZN(new_n146_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n147_));
  XNOR2_X1  g010(.A(new_n147_), .B(KEYINPUT2), .ZN(new_n148_));
  NAND2_X1  g011(.A1(new_n146_), .A2(new_n148_), .ZN(new_n149_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n150_));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n151_));
  INV_X1    g014(.A(new_n151_), .ZN(new_n152_));
  AND3_X1   g015(.A1(new_n149_), .A2(new_n150_), .A3(new_n152_), .ZN(new_n153_));
  AOI21_X1  g016(.A(new_n151_), .B1(KEYINPUT1), .B2(new_n150_), .ZN(new_n154_));
  OAI21_X1  g017(.A(new_n154_), .B1(KEYINPUT1), .B2(new_n150_), .ZN(new_n155_));
  INV_X1    g018(.A(new_n145_), .ZN(new_n156_));
  NAND3_X1  g019(.A1(new_n155_), .A2(new_n147_), .A3(new_n156_), .ZN(new_n157_));
  INV_X1    g020(.A(new_n157_), .ZN(new_n158_));
  OAI21_X1  g021(.A(new_n144_), .B1(new_n153_), .B2(new_n158_), .ZN(new_n159_));
  NAND3_X1  g022(.A1(new_n149_), .A2(new_n150_), .A3(new_n152_), .ZN(new_n160_));
  NAND4_X1  g023(.A1(new_n160_), .A2(new_n140_), .A3(new_n143_), .A4(new_n157_), .ZN(new_n161_));
  NAND3_X1  g024(.A1(new_n159_), .A2(KEYINPUT4), .A3(new_n161_), .ZN(new_n162_));
  NAND2_X1  g025(.A1(G225gat), .A2(G233gat), .ZN(new_n163_));
  INV_X1    g026(.A(new_n163_), .ZN(new_n164_));
  OAI211_X1 g027(.A(new_n162_), .B(new_n164_), .C1(KEYINPUT4), .C2(new_n159_), .ZN(new_n165_));
  NAND3_X1  g028(.A1(new_n159_), .A2(new_n163_), .A3(new_n161_), .ZN(new_n166_));
  NAND2_X1  g029(.A1(new_n165_), .A2(new_n166_), .ZN(new_n167_));
  XNOR2_X1  g030(.A(G1gat), .B(G29gat), .ZN(new_n168_));
  XNOR2_X1  g031(.A(new_n168_), .B(KEYINPUT0), .ZN(new_n169_));
  INV_X1    g032(.A(G57gat), .ZN(new_n170_));
  XNOR2_X1  g033(.A(new_n169_), .B(new_n170_), .ZN(new_n171_));
  INV_X1    g034(.A(G85gat), .ZN(new_n172_));
  XNOR2_X1  g035(.A(new_n171_), .B(new_n172_), .ZN(new_n173_));
  NAND2_X1  g036(.A1(new_n167_), .A2(new_n173_), .ZN(new_n174_));
  INV_X1    g037(.A(new_n173_), .ZN(new_n175_));
  NAND3_X1  g038(.A1(new_n175_), .A2(new_n165_), .A3(new_n166_), .ZN(new_n176_));
  NAND2_X1  g039(.A1(new_n174_), .A2(new_n176_), .ZN(new_n177_));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n178_));
  XNOR2_X1  g041(.A(new_n178_), .B(KEYINPUT23), .ZN(new_n179_));
  OAI21_X1  g042(.A(new_n179_), .B1(G183gat), .B2(G190gat), .ZN(new_n180_));
  INV_X1    g043(.A(G169gat), .ZN(new_n181_));
  INV_X1    g044(.A(G176gat), .ZN(new_n182_));
  NOR2_X1   g045(.A1(new_n181_), .A2(new_n182_), .ZN(new_n183_));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G169gat), .ZN(new_n184_));
  AOI21_X1  g047(.A(new_n183_), .B1(new_n184_), .B2(new_n182_), .ZN(new_n185_));
  NAND2_X1  g048(.A1(new_n180_), .A2(new_n185_), .ZN(new_n186_));
  XNOR2_X1  g049(.A(KEYINPUT25), .B(G183gat), .ZN(new_n187_));
  XNOR2_X1  g050(.A(KEYINPUT26), .B(G190gat), .ZN(new_n188_));
  NAND2_X1  g051(.A1(new_n187_), .A2(new_n188_), .ZN(new_n189_));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n190_));
  AOI21_X1  g053(.A(new_n190_), .B1(G169gat), .B2(G176gat), .ZN(new_n191_));
  OAI21_X1  g054(.A(new_n191_), .B1(G169gat), .B2(G176gat), .ZN(new_n192_));
  NAND3_X1  g055(.A1(new_n190_), .A2(new_n181_), .A3(new_n182_), .ZN(new_n193_));
  NAND4_X1  g056(.A1(new_n189_), .A2(new_n192_), .A3(new_n179_), .A4(new_n193_), .ZN(new_n194_));
  NAND2_X1  g057(.A1(new_n186_), .A2(new_n194_), .ZN(new_n195_));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n196_));
  XOR2_X1   g059(.A(G211gat), .B(G218gat), .Z(new_n197_));
  INV_X1    g060(.A(KEYINPUT21), .ZN(new_n198_));
  AOI21_X1  g061(.A(new_n196_), .B1(new_n197_), .B2(new_n198_), .ZN(new_n199_));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n200_));
  NAND2_X1  g063(.A1(new_n200_), .A2(KEYINPUT21), .ZN(new_n201_));
  NAND2_X1  g064(.A1(new_n199_), .A2(new_n201_), .ZN(new_n202_));
  NAND3_X1  g065(.A1(new_n200_), .A2(new_n196_), .A3(KEYINPUT21), .ZN(new_n203_));
  NAND2_X1  g066(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  AND2_X1   g067(.A1(new_n195_), .A2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g068(.A(KEYINPUT20), .B1(new_n195_), .B2(new_n204_), .ZN(new_n206_));
  NOR2_X1   g069(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XOR2_X1   g071(.A(new_n208_), .B(KEYINPUT19), .Z(new_n209_));
  NAND2_X1  g072(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g073(.A(new_n209_), .ZN(new_n211_));
  OAI21_X1  g074(.A(new_n211_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n212_));
  NAND2_X1  g075(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g076(.A(G8gat), .B(G36gat), .ZN(new_n214_));
  XNOR2_X1  g077(.A(new_n214_), .B(KEYINPUT18), .ZN(new_n215_));
  XNOR2_X1  g078(.A(new_n215_), .B(G64gat), .ZN(new_n216_));
  INV_X1    g079(.A(G92gat), .ZN(new_n217_));
  XNOR2_X1  g080(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  NAND3_X1  g081(.A1(new_n213_), .A2(KEYINPUT32), .A3(new_n218_), .ZN(new_n219_));
  AND2_X1   g082(.A1(new_n210_), .A2(new_n212_), .ZN(new_n220_));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n221_));
  INV_X1    g084(.A(new_n218_), .ZN(new_n222_));
  OAI21_X1  g085(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g086(.A1(new_n177_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n225_));
  NAND2_X1  g088(.A1(new_n176_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g089(.A1(new_n220_), .A2(new_n218_), .ZN(new_n227_));
  AOI21_X1  g090(.A(new_n218_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n228_));
  INV_X1    g091(.A(new_n228_), .ZN(new_n229_));
  OAI211_X1 g092(.A(new_n162_), .B(new_n163_), .C1(KEYINPUT4), .C2(new_n159_), .ZN(new_n230_));
  NAND3_X1  g093(.A1(new_n159_), .A2(new_n164_), .A3(new_n161_), .ZN(new_n231_));
  NAND3_X1  g094(.A1(new_n230_), .A2(new_n231_), .A3(new_n173_), .ZN(new_n232_));
  NAND4_X1  g095(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .A4(new_n232_), .ZN(new_n233_));
  NOR2_X1   g096(.A1(new_n176_), .A2(new_n225_), .ZN(new_n234_));
  OAI21_X1  g097(.A(new_n224_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n236_));
  XNOR2_X1  g099(.A(new_n236_), .B(KEYINPUT28), .ZN(new_n237_));
  XNOR2_X1  g100(.A(new_n237_), .B(G22gat), .ZN(new_n238_));
  AND2_X1   g101(.A1(new_n202_), .A2(new_n203_), .ZN(new_n239_));
  NAND2_X1  g102(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n240_));
  NOR2_X1   g103(.A1(new_n153_), .A2(new_n158_), .ZN(new_n241_));
  INV_X1    g104(.A(G228gat), .ZN(new_n242_));
  INV_X1    g105(.A(G233gat), .ZN(new_n243_));
  NOR2_X1   g106(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g107(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g108(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g109(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g110(.A(new_n245_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n248_));
  OAI21_X1  g111(.A(new_n238_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OR2_X1    g112(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n250_));
  INV_X1    g113(.A(G50gat), .ZN(new_n251_));
  XNOR2_X1  g114(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g115(.A1(new_n240_), .A2(new_n241_), .ZN(new_n253_));
  NAND2_X1  g116(.A1(new_n253_), .A2(new_n244_), .ZN(new_n254_));
  INV_X1    g117(.A(new_n238_), .ZN(new_n255_));
  NAND3_X1  g118(.A1(new_n254_), .A2(new_n246_), .A3(new_n255_), .ZN(new_n256_));
  AND3_X1   g119(.A1(new_n249_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g120(.A(new_n252_), .B1(new_n249_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g121(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g122(.A(G99gat), .ZN(new_n260_));
  XNOR2_X1  g123(.A(new_n144_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g124(.A(G15gat), .B(G43gat), .ZN(new_n262_));
  INV_X1    g125(.A(G71gat), .ZN(new_n263_));
  XNOR2_X1  g126(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  OR2_X1    g127(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g128(.A1(new_n261_), .A2(new_n264_), .ZN(new_n266_));
  NAND3_X1  g129(.A1(new_n265_), .A2(new_n195_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g130(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n269_));
  XOR2_X1   g132(.A(new_n269_), .B(KEYINPUT30), .Z(new_n270_));
  XNOR2_X1  g133(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  INV_X1    g134(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g135(.A(new_n195_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n273_));
  NOR3_X1   g136(.A1(new_n268_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g137(.A1(new_n265_), .A2(new_n266_), .ZN(new_n275_));
  INV_X1    g138(.A(new_n195_), .ZN(new_n276_));
  NAND2_X1  g139(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g140(.A(new_n271_), .B1(new_n277_), .B2(new_n267_), .ZN(new_n278_));
  NOR2_X1   g141(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g142(.A1(new_n259_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g143(.A1(new_n277_), .A2(new_n271_), .A3(new_n267_), .ZN(new_n281_));
  OAI21_X1  g144(.A(new_n272_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n282_));
  OAI211_X1 g145(.A(new_n281_), .B(new_n282_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n283_));
  INV_X1    g146(.A(new_n252_), .ZN(new_n284_));
  NOR3_X1   g147(.A1(new_n247_), .A2(new_n248_), .A3(new_n238_), .ZN(new_n285_));
  AOI21_X1  g148(.A(new_n255_), .B1(new_n254_), .B2(new_n246_), .ZN(new_n286_));
  OAI21_X1  g149(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g150(.A1(new_n249_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n288_));
  OAI211_X1 g151(.A(new_n287_), .B(new_n288_), .C1(new_n274_), .C2(new_n278_), .ZN(new_n289_));
  NAND2_X1  g152(.A1(new_n283_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g153(.A(KEYINPUT27), .ZN(new_n291_));
  NAND3_X1  g154(.A1(new_n227_), .A2(new_n229_), .A3(new_n291_), .ZN(new_n292_));
  NOR2_X1   g155(.A1(new_n213_), .A2(new_n222_), .ZN(new_n293_));
  OAI21_X1  g156(.A(KEYINPUT27), .B1(new_n293_), .B2(new_n228_), .ZN(new_n294_));
  AOI21_X1  g157(.A(new_n177_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g158(.A1(new_n235_), .A2(new_n280_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g159(.A(G15gat), .B(G22gat), .ZN(new_n297_));
  INV_X1    g160(.A(G1gat), .ZN(new_n298_));
  INV_X1    g161(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g162(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g163(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g164(.A(G1gat), .B(G8gat), .Z(new_n302_));
  XNOR2_X1  g165(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g166(.A(G43gat), .B(G50gat), .ZN(new_n304_));
  XNOR2_X1  g167(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g168(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g169(.A(new_n303_), .B(new_n306_), .ZN(new_n307_));
  NAND3_X1  g170(.A1(new_n307_), .A2(G229gat), .A3(G233gat), .ZN(new_n308_));
  NAND2_X1  g171(.A1(G229gat), .A2(G233gat), .ZN(new_n309_));
  NAND2_X1  g172(.A1(new_n303_), .A2(new_n306_), .ZN(new_n310_));
  INV_X1    g173(.A(KEYINPUT15), .ZN(new_n311_));
  XNOR2_X1  g174(.A(new_n306_), .B(new_n311_), .ZN(new_n312_));
  OAI211_X1 g175(.A(new_n309_), .B(new_n310_), .C1(new_n312_), .C2(new_n303_), .ZN(new_n313_));
  NAND2_X1  g176(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g177(.A(G113gat), .B(G141gat), .ZN(new_n315_));
  XNOR2_X1  g178(.A(G169gat), .B(G197gat), .ZN(new_n316_));
  XOR2_X1   g179(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  INV_X1    g180(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g181(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g182(.A1(new_n308_), .A2(new_n317_), .A3(new_n313_), .ZN(new_n320_));
  NAND2_X1  g183(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g184(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g185(.A(KEYINPUT36), .ZN(new_n323_));
  XNOR2_X1  g186(.A(G85gat), .B(G92gat), .ZN(new_n324_));
  INV_X1    g187(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g188(.A1(G99gat), .A2(G106gat), .ZN(new_n326_));
  NAND2_X1  g189(.A1(new_n326_), .A2(KEYINPUT6), .ZN(new_n327_));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n328_));
  NAND3_X1  g191(.A1(new_n328_), .A2(G99gat), .A3(G106gat), .ZN(new_n329_));
  AND2_X1   g192(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g193(.A(KEYINPUT7), .ZN(new_n331_));
  INV_X1    g194(.A(G106gat), .ZN(new_n332_));
  NAND3_X1  g195(.A1(new_n331_), .A2(new_n260_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g196(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n334_));
  NAND2_X1  g197(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g198(.A(new_n325_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g199(.A1(new_n336_), .A2(KEYINPUT8), .ZN(new_n337_));
  AOI21_X1  g200(.A(new_n328_), .B1(G99gat), .B2(G106gat), .ZN(new_n338_));
  NOR2_X1   g201(.A1(new_n326_), .A2(KEYINPUT6), .ZN(new_n339_));
  OAI211_X1 g202(.A(new_n334_), .B(new_n333_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g203(.A(KEYINPUT8), .ZN(new_n341_));
  NAND3_X1  g204(.A1(new_n340_), .A2(new_n341_), .A3(new_n325_), .ZN(new_n342_));
  NAND2_X1  g205(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g206(.A(KEYINPUT10), .B(G99gat), .ZN(new_n344_));
  OR2_X1    g207(.A1(new_n344_), .A2(G106gat), .ZN(new_n345_));
  NAND2_X1  g208(.A1(new_n327_), .A2(new_n329_), .ZN(new_n346_));
  INV_X1    g209(.A(KEYINPUT9), .ZN(new_n347_));
  OAI21_X1  g210(.A(new_n347_), .B1(new_n172_), .B2(new_n217_), .ZN(new_n348_));
  NAND3_X1  g211(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n349_));
  OAI211_X1 g212(.A(new_n348_), .B(new_n349_), .C1(G85gat), .C2(G92gat), .ZN(new_n350_));
  NAND3_X1  g213(.A1(new_n345_), .A2(new_n346_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g214(.A1(new_n343_), .A2(new_n306_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g215(.A1(G232gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g216(.A(new_n353_), .B(KEYINPUT34), .Z(new_n354_));
  INV_X1    g217(.A(KEYINPUT35), .ZN(new_n355_));
  NAND2_X1  g218(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g219(.A1(new_n345_), .A2(new_n350_), .A3(new_n346_), .ZN(new_n357_));
  AOI21_X1  g220(.A(new_n357_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n358_));
  OAI211_X1 g221(.A(new_n352_), .B(new_n356_), .C1(new_n312_), .C2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g222(.A1(new_n354_), .A2(new_n355_), .ZN(new_n360_));
  NOR2_X1   g223(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g224(.A(new_n360_), .ZN(new_n362_));
  XNOR2_X1  g225(.A(new_n306_), .B(KEYINPUT15), .ZN(new_n363_));
  INV_X1    g226(.A(new_n334_), .ZN(new_n364_));
  NOR3_X1   g227(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n365_));
  NOR2_X1   g228(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI211_X1 g229(.A(KEYINPUT8), .B(new_n324_), .C1(new_n366_), .C2(new_n346_), .ZN(new_n367_));
  AOI21_X1  g230(.A(new_n341_), .B1(new_n340_), .B2(new_n325_), .ZN(new_n368_));
  OAI21_X1  g231(.A(new_n351_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g232(.A1(new_n363_), .A2(new_n369_), .B1(new_n355_), .B2(new_n354_), .ZN(new_n370_));
  AOI21_X1  g233(.A(new_n362_), .B1(new_n370_), .B2(new_n352_), .ZN(new_n371_));
  OAI21_X1  g234(.A(new_n323_), .B1(new_n361_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g235(.A(G134gat), .B(G162gat), .ZN(new_n373_));
  XNOR2_X1  g236(.A(new_n373_), .B(G190gat), .ZN(new_n374_));
  XNOR2_X1  g237(.A(new_n374_), .B(G218gat), .ZN(new_n375_));
  INV_X1    g238(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g239(.A1(new_n359_), .A2(new_n360_), .ZN(new_n377_));
  NAND3_X1  g240(.A1(new_n370_), .A2(new_n352_), .A3(new_n362_), .ZN(new_n378_));
  NAND3_X1  g241(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT36), .ZN(new_n379_));
  NAND3_X1  g242(.A1(new_n372_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  OAI211_X1 g243(.A(new_n323_), .B(new_n375_), .C1(new_n361_), .C2(new_n371_), .ZN(new_n381_));
  NAND2_X1  g244(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n383_));
  NAND2_X1  g246(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g247(.A(G78gat), .ZN(new_n385_));
  NAND2_X1  g248(.A1(new_n263_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g249(.A1(G71gat), .A2(G78gat), .ZN(new_n387_));
  NAND2_X1  g250(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n389_));
  NAND2_X1  g252(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g253(.A1(new_n386_), .A2(KEYINPUT11), .A3(new_n387_), .ZN(new_n391_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n392_));
  NAND3_X1  g255(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  OR2_X1    g256(.A1(new_n391_), .A2(new_n392_), .ZN(new_n394_));
  NAND2_X1  g257(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g258(.A(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g259(.A(new_n396_), .B(new_n303_), .ZN(new_n397_));
  NAND2_X1  g260(.A1(G231gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g261(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g262(.A(G183gat), .B(G211gat), .ZN(new_n400_));
  XNOR2_X1  g263(.A(new_n400_), .B(KEYINPUT16), .ZN(new_n401_));
  XNOR2_X1  g264(.A(G127gat), .B(G155gat), .ZN(new_n402_));
  XNOR2_X1  g265(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g266(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n405_));
  NAND2_X1  g268(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g269(.A1(new_n399_), .A2(KEYINPUT17), .A3(new_n403_), .ZN(new_n407_));
  OR2_X1    g270(.A1(new_n399_), .A2(new_n403_), .ZN(new_n408_));
  NAND3_X1  g271(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g272(.A1(new_n380_), .A2(KEYINPUT37), .A3(new_n381_), .ZN(new_n410_));
  NAND3_X1  g273(.A1(new_n384_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NOR3_X1   g274(.A1(new_n296_), .A2(new_n322_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g275(.A1(G230gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g276(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g277(.A1(new_n369_), .A2(new_n396_), .ZN(new_n415_));
  OAI211_X1 g278(.A(new_n351_), .B(new_n395_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n416_));
  NAND3_X1  g279(.A1(new_n415_), .A2(KEYINPUT12), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n418_));
  NAND3_X1  g281(.A1(new_n369_), .A2(new_n418_), .A3(new_n396_), .ZN(new_n419_));
  AOI21_X1  g282(.A(new_n414_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g283(.A(G176gat), .B(G204gat), .ZN(new_n421_));
  XNOR2_X1  g284(.A(new_n421_), .B(KEYINPUT5), .ZN(new_n422_));
  XNOR2_X1  g285(.A(new_n422_), .B(G120gat), .ZN(new_n423_));
  XOR2_X1   g286(.A(new_n423_), .B(G148gat), .Z(new_n424_));
  AOI21_X1  g287(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n425_));
  NOR3_X1   g288(.A1(new_n420_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g289(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g290(.A(new_n424_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n428_));
  NAND3_X1  g291(.A1(new_n427_), .A2(KEYINPUT13), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n430_));
  INV_X1    g293(.A(new_n428_), .ZN(new_n431_));
  OAI21_X1  g294(.A(new_n430_), .B1(new_n431_), .B2(new_n426_), .ZN(new_n432_));
  NAND2_X1  g295(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g296(.A(new_n177_), .ZN(new_n434_));
  NOR2_X1   g297(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g298(.A1(new_n412_), .A2(new_n298_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g299(.A(new_n436_), .B(KEYINPUT38), .ZN(new_n437_));
  INV_X1    g300(.A(new_n382_), .ZN(new_n438_));
  INV_X1    g301(.A(new_n409_), .ZN(new_n439_));
  NOR3_X1   g302(.A1(new_n296_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g303(.A1(new_n433_), .A2(new_n322_), .ZN(new_n441_));
  NAND2_X1  g304(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g305(.A(G1gat), .B1(new_n442_), .B2(new_n434_), .ZN(new_n443_));
  NAND2_X1  g306(.A1(new_n437_), .A2(new_n443_), .ZN(G1324gat));
  NAND2_X1  g307(.A1(new_n292_), .A2(new_n294_), .ZN(new_n445_));
  NOR2_X1   g308(.A1(new_n433_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g309(.A1(new_n412_), .A2(new_n299_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g310(.A(G8gat), .B1(new_n442_), .B2(new_n445_), .ZN(new_n448_));
  AND2_X1   g311(.A1(new_n448_), .A2(KEYINPUT39), .ZN(new_n449_));
  NOR2_X1   g312(.A1(new_n448_), .A2(KEYINPUT39), .ZN(new_n450_));
  OAI21_X1  g313(.A(new_n447_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n452_));
  NAND2_X1  g315(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g316(.A(KEYINPUT40), .B(new_n447_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n454_));
  NAND2_X1  g317(.A1(new_n453_), .A2(new_n454_), .ZN(G1325gat));
  INV_X1    g318(.A(new_n279_), .ZN(new_n456_));
  OAI21_X1  g319(.A(G15gat), .B1(new_n442_), .B2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g320(.A(new_n457_), .B(KEYINPUT41), .Z(new_n458_));
  INV_X1    g321(.A(G15gat), .ZN(new_n459_));
  NOR2_X1   g322(.A1(new_n433_), .A2(new_n456_), .ZN(new_n460_));
  NAND3_X1  g323(.A1(new_n412_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g324(.A1(new_n458_), .A2(new_n461_), .ZN(G1326gat));
  INV_X1    g325(.A(new_n259_), .ZN(new_n463_));
  OAI21_X1  g326(.A(G22gat), .B1(new_n442_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g327(.A(new_n464_), .B(KEYINPUT42), .ZN(new_n465_));
  INV_X1    g328(.A(G22gat), .ZN(new_n466_));
  NOR2_X1   g329(.A1(new_n433_), .A2(new_n463_), .ZN(new_n467_));
  NAND3_X1  g330(.A1(new_n412_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g331(.A1(new_n465_), .A2(new_n468_), .ZN(G1327gat));
  NOR2_X1   g332(.A1(new_n296_), .A2(new_n322_), .ZN(new_n470_));
  NOR2_X1   g333(.A1(new_n409_), .A2(new_n382_), .ZN(new_n471_));
  NAND2_X1  g334(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g335(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g336(.A(G29gat), .ZN(new_n474_));
  NAND3_X1  g337(.A1(new_n473_), .A2(new_n474_), .A3(new_n435_), .ZN(new_n475_));
  INV_X1    g338(.A(new_n410_), .ZN(new_n476_));
  AOI21_X1  g339(.A(KEYINPUT37), .B1(new_n380_), .B2(new_n381_), .ZN(new_n477_));
  NOR2_X1   g340(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g341(.A(KEYINPUT43), .B1(new_n296_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g342(.A1(new_n235_), .A2(new_n280_), .ZN(new_n480_));
  NAND2_X1  g343(.A1(new_n290_), .A2(new_n295_), .ZN(new_n481_));
  NAND2_X1  g344(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g345(.A(KEYINPUT43), .ZN(new_n483_));
  NAND2_X1  g346(.A1(new_n384_), .A2(new_n410_), .ZN(new_n484_));
  NAND3_X1  g347(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g348(.A1(new_n479_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g349(.A1(new_n441_), .A2(new_n439_), .ZN(new_n487_));
  INV_X1    g350(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g351(.A(KEYINPUT44), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g352(.A(KEYINPUT44), .ZN(new_n490_));
  AOI211_X1 g353(.A(new_n490_), .B(new_n487_), .C1(new_n479_), .C2(new_n485_), .ZN(new_n491_));
  NOR3_X1   g354(.A1(new_n489_), .A2(new_n491_), .A3(new_n434_), .ZN(new_n492_));
  OAI21_X1  g355(.A(new_n475_), .B1(new_n492_), .B2(new_n474_), .ZN(G1328gat));
  INV_X1    g356(.A(KEYINPUT46), .ZN(new_n494_));
  INV_X1    g357(.A(G36gat), .ZN(new_n495_));
  NOR2_X1   g358(.A1(new_n489_), .A2(new_n491_), .ZN(new_n496_));
  INV_X1    g359(.A(new_n445_), .ZN(new_n497_));
  AOI21_X1  g360(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g361(.A1(new_n446_), .A2(new_n495_), .ZN(new_n499_));
  OR3_X1    g362(.A1(new_n472_), .A2(KEYINPUT45), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g363(.A(KEYINPUT45), .B1(new_n472_), .B2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g364(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g365(.A(new_n502_), .ZN(new_n503_));
  OAI21_X1  g366(.A(new_n494_), .B1(new_n498_), .B2(new_n503_), .ZN(new_n504_));
  NOR3_X1   g367(.A1(new_n489_), .A2(new_n491_), .A3(new_n445_), .ZN(new_n505_));
  OAI211_X1 g368(.A(KEYINPUT46), .B(new_n502_), .C1(new_n505_), .C2(new_n495_), .ZN(new_n506_));
  NAND2_X1  g369(.A1(new_n504_), .A2(new_n506_), .ZN(G1329gat));
  INV_X1    g370(.A(KEYINPUT47), .ZN(new_n508_));
  INV_X1    g371(.A(G43gat), .ZN(new_n509_));
  AOI21_X1  g372(.A(new_n509_), .B1(new_n496_), .B2(new_n279_), .ZN(new_n510_));
  NAND2_X1  g373(.A1(new_n460_), .A2(new_n509_), .ZN(new_n511_));
  NOR2_X1   g374(.A1(new_n472_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g375(.A(new_n508_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NOR3_X1   g376(.A1(new_n489_), .A2(new_n491_), .A3(new_n456_), .ZN(new_n514_));
  OAI221_X1 g377(.A(KEYINPUT47), .B1(new_n472_), .B2(new_n511_), .C1(new_n514_), .C2(new_n509_), .ZN(new_n515_));
  NAND2_X1  g378(.A1(new_n513_), .A2(new_n515_), .ZN(G1330gat));
  NAND3_X1  g379(.A1(new_n473_), .A2(new_n251_), .A3(new_n467_), .ZN(new_n517_));
  NOR3_X1   g380(.A1(new_n489_), .A2(new_n491_), .A3(new_n463_), .ZN(new_n518_));
  OAI21_X1  g381(.A(new_n517_), .B1(new_n518_), .B2(new_n251_), .ZN(G1331gat));
  NOR3_X1   g382(.A1(new_n296_), .A2(new_n321_), .A3(new_n411_), .ZN(new_n520_));
  INV_X1    g383(.A(new_n433_), .ZN(new_n521_));
  NOR2_X1   g384(.A1(new_n521_), .A2(new_n434_), .ZN(new_n522_));
  NAND3_X1  g385(.A1(new_n520_), .A2(new_n170_), .A3(new_n522_), .ZN(new_n523_));
  NOR2_X1   g386(.A1(new_n521_), .A2(new_n321_), .ZN(new_n524_));
  AND2_X1   g387(.A1(new_n440_), .A2(new_n524_), .ZN(new_n525_));
  AND2_X1   g388(.A1(new_n525_), .A2(new_n177_), .ZN(new_n526_));
  OAI21_X1  g389(.A(new_n523_), .B1(new_n526_), .B2(new_n170_), .ZN(G1332gat));
  INV_X1    g390(.A(G64gat), .ZN(new_n528_));
  AOI21_X1  g391(.A(new_n528_), .B1(new_n525_), .B2(new_n497_), .ZN(new_n529_));
  XOR2_X1   g392(.A(new_n529_), .B(KEYINPUT48), .Z(new_n530_));
  NOR2_X1   g393(.A1(new_n521_), .A2(new_n445_), .ZN(new_n531_));
  NAND3_X1  g394(.A1(new_n520_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g395(.A1(new_n530_), .A2(new_n532_), .ZN(G1333gat));
  AOI21_X1  g396(.A(new_n263_), .B1(new_n525_), .B2(new_n279_), .ZN(new_n534_));
  XOR2_X1   g397(.A(new_n534_), .B(KEYINPUT49), .Z(new_n535_));
  NOR2_X1   g398(.A1(new_n521_), .A2(new_n456_), .ZN(new_n536_));
  NAND3_X1  g399(.A1(new_n520_), .A2(new_n263_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g400(.A1(new_n535_), .A2(new_n537_), .ZN(G1334gat));
  AOI21_X1  g401(.A(new_n385_), .B1(new_n525_), .B2(new_n259_), .ZN(new_n539_));
  XOR2_X1   g402(.A(new_n539_), .B(KEYINPUT50), .Z(new_n540_));
  NOR2_X1   g403(.A1(new_n521_), .A2(new_n463_), .ZN(new_n541_));
  NAND3_X1  g404(.A1(new_n520_), .A2(new_n385_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g405(.A1(new_n540_), .A2(new_n542_), .ZN(G1335gat));
  NOR2_X1   g406(.A1(new_n296_), .A2(new_n321_), .ZN(new_n544_));
  NAND2_X1  g407(.A1(new_n544_), .A2(new_n471_), .ZN(new_n545_));
  INV_X1    g408(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g409(.A1(new_n546_), .A2(new_n172_), .A3(new_n522_), .ZN(new_n547_));
  AND3_X1   g410(.A1(new_n486_), .A2(new_n439_), .A3(new_n524_), .ZN(new_n548_));
  AND2_X1   g411(.A1(new_n548_), .A2(new_n177_), .ZN(new_n549_));
  OAI21_X1  g412(.A(new_n547_), .B1(new_n549_), .B2(new_n172_), .ZN(G1336gat));
  NAND3_X1  g413(.A1(new_n546_), .A2(new_n217_), .A3(new_n531_), .ZN(new_n551_));
  AND2_X1   g414(.A1(new_n548_), .A2(new_n497_), .ZN(new_n552_));
  OAI21_X1  g415(.A(new_n551_), .B1(new_n552_), .B2(new_n217_), .ZN(G1337gat));
  AOI21_X1  g416(.A(new_n260_), .B1(new_n548_), .B2(new_n279_), .ZN(new_n554_));
  NOR4_X1   g417(.A1(new_n545_), .A2(new_n344_), .A3(new_n521_), .A4(new_n456_), .ZN(new_n555_));
  OR3_X1    g418(.A1(new_n554_), .A2(KEYINPUT51), .A3(new_n555_), .ZN(new_n556_));
  OAI21_X1  g419(.A(KEYINPUT51), .B1(new_n554_), .B2(new_n555_), .ZN(new_n557_));
  NAND2_X1  g420(.A1(new_n556_), .A2(new_n557_), .ZN(G1338gat));
  NAND3_X1  g421(.A1(new_n546_), .A2(new_n332_), .A3(new_n541_), .ZN(new_n559_));
  NAND4_X1  g422(.A1(new_n486_), .A2(new_n259_), .A3(new_n439_), .A4(new_n524_), .ZN(new_n560_));
  INV_X1    g423(.A(KEYINPUT52), .ZN(new_n561_));
  AND3_X1   g424(.A1(new_n560_), .A2(new_n561_), .A3(G106gat), .ZN(new_n562_));
  AOI21_X1  g425(.A(new_n561_), .B1(new_n560_), .B2(G106gat), .ZN(new_n563_));
  OAI21_X1  g426(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g427(.A1(new_n564_), .A2(KEYINPUT53), .ZN(new_n565_));
  INV_X1    g428(.A(KEYINPUT53), .ZN(new_n566_));
  OAI211_X1 g429(.A(new_n566_), .B(new_n559_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g430(.A1(new_n565_), .A2(new_n567_), .ZN(G1339gat));
  NAND3_X1  g431(.A1(new_n429_), .A2(new_n432_), .A3(new_n322_), .ZN(new_n569_));
  OAI21_X1  g432(.A(KEYINPUT54), .B1(new_n411_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g433(.A(new_n569_), .ZN(new_n571_));
  INV_X1    g434(.A(KEYINPUT54), .ZN(new_n572_));
  NAND4_X1  g435(.A1(new_n478_), .A2(new_n571_), .A3(new_n572_), .A4(new_n409_), .ZN(new_n573_));
  AND2_X1   g436(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g437(.A1(new_n427_), .A2(new_n321_), .ZN(new_n575_));
  INV_X1    g438(.A(KEYINPUT56), .ZN(new_n576_));
  NAND3_X1  g439(.A1(new_n417_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n577_));
  INV_X1    g440(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g441(.A1(new_n416_), .A2(KEYINPUT12), .ZN(new_n579_));
  AOI21_X1  g442(.A(new_n395_), .B1(new_n343_), .B2(new_n351_), .ZN(new_n580_));
  NOR2_X1   g443(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g444(.A(new_n419_), .ZN(new_n582_));
  OAI21_X1  g445(.A(new_n413_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g446(.A1(new_n583_), .A2(KEYINPUT55), .ZN(new_n584_));
  INV_X1    g447(.A(KEYINPUT55), .ZN(new_n585_));
  NAND2_X1  g448(.A1(new_n420_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g449(.A(new_n578_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g450(.A(new_n424_), .ZN(new_n588_));
  OAI21_X1  g451(.A(new_n576_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g452(.A1(new_n417_), .A2(new_n419_), .ZN(new_n590_));
  AOI21_X1  g453(.A(new_n585_), .B1(new_n590_), .B2(new_n413_), .ZN(new_n591_));
  AOI211_X1 g454(.A(KEYINPUT55), .B(new_n414_), .C1(new_n417_), .C2(new_n419_), .ZN(new_n592_));
  OAI21_X1  g455(.A(new_n577_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g456(.A1(new_n593_), .A2(KEYINPUT56), .A3(new_n424_), .ZN(new_n594_));
  AOI21_X1  g457(.A(new_n575_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g458(.A(new_n317_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n596_));
  OAI21_X1  g459(.A(new_n310_), .B1(new_n312_), .B2(new_n303_), .ZN(new_n597_));
  OAI21_X1  g460(.A(new_n596_), .B1(new_n309_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g461(.A1(new_n598_), .A2(new_n320_), .ZN(new_n599_));
  AOI21_X1  g462(.A(new_n599_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n600_));
  OAI21_X1  g463(.A(new_n382_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g464(.A(KEYINPUT57), .ZN(new_n602_));
  NAND2_X1  g465(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g466(.A1(new_n426_), .A2(new_n599_), .ZN(new_n604_));
  AND3_X1   g467(.A1(new_n593_), .A2(KEYINPUT56), .A3(new_n424_), .ZN(new_n605_));
  AOI21_X1  g468(.A(KEYINPUT56), .B1(new_n593_), .B2(new_n424_), .ZN(new_n606_));
  OAI21_X1  g469(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g470(.A(KEYINPUT58), .ZN(new_n608_));
  NAND2_X1  g471(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g472(.A(KEYINPUT58), .B(new_n604_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n610_));
  NAND3_X1  g473(.A1(new_n609_), .A2(new_n484_), .A3(new_n610_), .ZN(new_n611_));
  OAI211_X1 g474(.A(KEYINPUT57), .B(new_n382_), .C1(new_n595_), .C2(new_n600_), .ZN(new_n612_));
  NAND3_X1  g475(.A1(new_n603_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g476(.A(new_n574_), .B1(new_n613_), .B2(new_n439_), .ZN(new_n614_));
  NOR2_X1   g477(.A1(new_n497_), .A2(new_n283_), .ZN(new_n615_));
  INV_X1    g478(.A(new_n615_), .ZN(new_n616_));
  NOR3_X1   g479(.A1(new_n614_), .A2(new_n434_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g480(.A(G113gat), .ZN(new_n618_));
  NAND3_X1  g481(.A1(new_n617_), .A2(new_n618_), .A3(new_n321_), .ZN(new_n619_));
  INV_X1    g482(.A(KEYINPUT59), .ZN(new_n620_));
  NAND2_X1  g483(.A1(new_n613_), .A2(new_n439_), .ZN(new_n621_));
  INV_X1    g484(.A(new_n574_), .ZN(new_n622_));
  AOI21_X1  g485(.A(new_n434_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g486(.A(new_n620_), .B1(new_n623_), .B2(new_n615_), .ZN(new_n624_));
  NOR4_X1   g487(.A1(new_n614_), .A2(KEYINPUT59), .A3(new_n434_), .A4(new_n616_), .ZN(new_n625_));
  NOR3_X1   g488(.A1(new_n624_), .A2(new_n625_), .A3(new_n322_), .ZN(new_n626_));
  OAI21_X1  g489(.A(new_n619_), .B1(new_n626_), .B2(new_n618_), .ZN(G1340gat));
  INV_X1    g490(.A(G120gat), .ZN(new_n628_));
  AOI21_X1  g491(.A(KEYINPUT60), .B1(new_n433_), .B2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g492(.A(new_n629_), .B1(KEYINPUT60), .B2(new_n628_), .ZN(new_n630_));
  NAND2_X1  g493(.A1(new_n617_), .A2(new_n630_), .ZN(new_n631_));
  NOR3_X1   g494(.A1(new_n624_), .A2(new_n625_), .A3(new_n521_), .ZN(new_n632_));
  OAI21_X1  g495(.A(new_n631_), .B1(new_n632_), .B2(new_n628_), .ZN(G1341gat));
  INV_X1    g496(.A(G127gat), .ZN(new_n634_));
  NAND3_X1  g497(.A1(new_n617_), .A2(new_n634_), .A3(new_n409_), .ZN(new_n635_));
  NOR3_X1   g498(.A1(new_n624_), .A2(new_n625_), .A3(new_n439_), .ZN(new_n636_));
  OAI21_X1  g499(.A(new_n635_), .B1(new_n636_), .B2(new_n634_), .ZN(G1342gat));
  INV_X1    g500(.A(G134gat), .ZN(new_n638_));
  NAND3_X1  g501(.A1(new_n617_), .A2(new_n638_), .A3(new_n438_), .ZN(new_n639_));
  NOR3_X1   g502(.A1(new_n624_), .A2(new_n625_), .A3(new_n478_), .ZN(new_n640_));
  OAI21_X1  g503(.A(new_n639_), .B1(new_n640_), .B2(new_n638_), .ZN(G1343gat));
  NOR4_X1   g504(.A1(new_n614_), .A2(new_n434_), .A3(new_n289_), .A4(new_n497_), .ZN(new_n642_));
  NAND2_X1  g505(.A1(new_n642_), .A2(new_n321_), .ZN(new_n643_));
  XNOR2_X1  g506(.A(new_n643_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g507(.A1(new_n642_), .A2(new_n433_), .ZN(new_n645_));
  XNOR2_X1  g508(.A(new_n645_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g509(.A1(new_n642_), .A2(new_n409_), .ZN(new_n647_));
  XNOR2_X1  g510(.A(KEYINPUT61), .B(G155gat), .ZN(new_n648_));
  XNOR2_X1  g511(.A(new_n647_), .B(new_n648_), .ZN(G1346gat));
  INV_X1    g512(.A(G162gat), .ZN(new_n650_));
  NAND3_X1  g513(.A1(new_n642_), .A2(new_n650_), .A3(new_n438_), .ZN(new_n651_));
  AND2_X1   g514(.A1(new_n642_), .A2(new_n484_), .ZN(new_n652_));
  OAI21_X1  g515(.A(new_n651_), .B1(new_n652_), .B2(new_n650_), .ZN(G1347gat));
  AOI21_X1  g516(.A(new_n177_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n654_));
  INV_X1    g517(.A(new_n283_), .ZN(new_n655_));
  NAND4_X1  g518(.A1(new_n654_), .A2(new_n321_), .A3(new_n655_), .A4(new_n497_), .ZN(new_n656_));
  NAND2_X1  g519(.A1(new_n656_), .A2(G169gat), .ZN(new_n657_));
  INV_X1    g520(.A(KEYINPUT62), .ZN(new_n658_));
  NAND2_X1  g521(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g522(.A1(new_n656_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n660_));
  NOR3_X1   g523(.A1(new_n614_), .A2(new_n177_), .A3(new_n283_), .ZN(new_n661_));
  NAND4_X1  g524(.A1(new_n661_), .A2(new_n321_), .A3(new_n184_), .A4(new_n497_), .ZN(new_n662_));
  NAND3_X1  g525(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(G1348gat));
  NAND2_X1  g526(.A1(new_n661_), .A2(new_n531_), .ZN(new_n664_));
  XNOR2_X1  g527(.A(new_n664_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g528(.A1(new_n661_), .A2(new_n497_), .ZN(new_n666_));
  OAI21_X1  g529(.A(G183gat), .B1(new_n666_), .B2(new_n439_), .ZN(new_n667_));
  NAND4_X1  g530(.A1(new_n661_), .A2(new_n187_), .A3(new_n497_), .A4(new_n409_), .ZN(new_n668_));
  NAND2_X1  g531(.A1(new_n667_), .A2(new_n668_), .ZN(G1350gat));
  OAI21_X1  g532(.A(G190gat), .B1(new_n666_), .B2(new_n478_), .ZN(new_n670_));
  NAND2_X1  g533(.A1(new_n438_), .A2(new_n188_), .ZN(new_n671_));
  OAI21_X1  g534(.A(new_n670_), .B1(new_n666_), .B2(new_n671_), .ZN(G1351gat));
  NOR3_X1   g535(.A1(new_n614_), .A2(new_n177_), .A3(new_n289_), .ZN(new_n673_));
  NAND3_X1  g536(.A1(new_n673_), .A2(new_n321_), .A3(new_n497_), .ZN(new_n674_));
  XNOR2_X1  g537(.A(new_n674_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g538(.A1(new_n673_), .A2(new_n531_), .ZN(new_n676_));
  XNOR2_X1  g539(.A(new_n676_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g540(.A(new_n439_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n678_));
  NAND3_X1  g541(.A1(new_n673_), .A2(new_n497_), .A3(new_n678_), .ZN(new_n679_));
  OR2_X1    g542(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n680_));
  XNOR2_X1  g543(.A(new_n679_), .B(new_n680_), .ZN(G1354gat));
  NAND3_X1  g544(.A1(new_n673_), .A2(new_n497_), .A3(new_n484_), .ZN(new_n682_));
  NAND2_X1  g545(.A1(new_n682_), .A2(G218gat), .ZN(new_n683_));
  NOR2_X1   g546(.A1(new_n382_), .A2(G218gat), .ZN(new_n684_));
  NAND3_X1  g547(.A1(new_n673_), .A2(new_n497_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g548(.A1(new_n683_), .A2(new_n685_), .ZN(G1355gat));
endmodule


