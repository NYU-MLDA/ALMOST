//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n991_, new_n992_, new_n994_, new_n995_, new_n996_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1005_, new_n1006_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT19), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT25), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G190gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(KEYINPUT24), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT79), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT23), .ZN(new_n230_));
  AND2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n231_), .B2(new_n227_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n227_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(new_n231_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n210_), .A2(new_n214_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n219_), .A2(KEYINPUT22), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G169gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n245_), .A3(new_n220_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n246_), .A2(new_n222_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n226_), .A2(new_n237_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(G197gat), .A2(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT21), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G218gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G211gat), .ZN(new_n256_));
  INV_X1    g055(.A(G211gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G218gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n251_), .B(new_n254_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n254_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n256_), .A2(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT88), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n209_), .B1(new_n248_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n242_), .A2(new_n247_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n225_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n237_), .A2(new_n271_), .A3(new_n218_), .A4(new_n223_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n262_), .A2(new_n267_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(KEYINPUT90), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT78), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n218_), .A2(new_n278_), .A3(new_n223_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n228_), .A2(new_n230_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n235_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n225_), .B1(new_n281_), .B2(new_n238_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n237_), .A2(new_n241_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n246_), .A2(KEYINPUT80), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n246_), .A2(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n268_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(KEYINPUT20), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n208_), .B1(new_n276_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n248_), .B2(new_n268_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n283_), .A2(new_n287_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n292_), .B(new_n208_), .C1(new_n268_), .C2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n205_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G29gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(G85gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G57gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT84), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n305_));
  INV_X1    g104(.A(G134gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G127gat), .ZN(new_n307_));
  INV_X1    g106(.A(G127gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G134gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G120gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G113gat), .ZN(new_n312_));
  INV_X1    g111(.A(G113gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G120gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n305_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n304_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  INV_X1    g117(.A(G141gat), .ZN(new_n319_));
  INV_X1    g118(.A(G148gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n322_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(new_n339_), .A3(new_n329_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n335_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n331_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n307_), .A2(new_n309_), .A3(new_n312_), .A4(new_n314_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT83), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n302_), .A2(new_n303_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n317_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n337_), .B1(new_n334_), .B2(new_n333_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n349_), .A2(new_n340_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n310_), .A2(new_n315_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n307_), .A2(new_n309_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT91), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n310_), .A2(new_n315_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT91), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n343_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n348_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n348_), .A2(new_n357_), .A3(KEYINPUT4), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n317_), .A2(new_n342_), .A3(new_n361_), .A4(new_n347_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n301_), .B(new_n359_), .C1(new_n360_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT33), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n348_), .A2(new_n357_), .A3(KEYINPUT4), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(new_n363_), .A3(new_n362_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n301_), .A4(new_n359_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n205_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n288_), .A2(KEYINPUT20), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n372_), .B(new_n294_), .C1(new_n374_), .C2(new_n208_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n348_), .A2(new_n357_), .A3(new_n363_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n300_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n362_), .A2(new_n358_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n377_), .A2(new_n378_), .B1(new_n379_), .B2(new_n367_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(KEYINPUT92), .A3(new_n300_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n296_), .A2(new_n371_), .A3(new_n375_), .A4(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n365_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n301_), .B1(new_n368_), .B2(new_n359_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n372_), .A2(KEYINPUT32), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n294_), .B(new_n390_), .C1(new_n374_), .C2(new_n208_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n292_), .B1(new_n268_), .B2(new_n293_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n207_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n276_), .A2(new_n289_), .A3(new_n208_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n389_), .B(new_n391_), .C1(new_n390_), .C2(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n366_), .A2(new_n370_), .B1(new_n381_), .B2(new_n380_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n397_), .A2(KEYINPUT93), .A3(new_n375_), .A4(new_n296_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n385_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n400_), .B(new_n274_), .C1(new_n401_), .C2(KEYINPUT86), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n403_), .A2(KEYINPUT87), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n401_), .B(new_n274_), .C1(KEYINPUT86), .C2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n411_));
  XOR2_X1   g210(.A(G22gat), .B(G50gat), .Z(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT28), .Z(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n404_), .A2(new_n407_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n405_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n408_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n418_), .A2(KEYINPUT89), .A3(new_n408_), .A4(new_n414_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n375_), .A2(KEYINPUT27), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n372_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT27), .B1(new_n296_), .B2(new_n375_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n422_), .A2(new_n389_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n399_), .A2(new_n422_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT31), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n293_), .B(KEYINPUT30), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434_));
  INV_X1    g233(.A(G43gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(G15gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n436_), .B(new_n439_), .Z(new_n440_));
  AOI21_X1  g239(.A(new_n430_), .B1(new_n433_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n430_), .A3(new_n440_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n293_), .B(KEYINPUT30), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n317_), .A2(new_n347_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(KEYINPUT82), .A3(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n347_), .B(new_n317_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n442_), .A2(new_n443_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n447_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n443_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n441_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n427_), .A2(new_n422_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n388_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n429_), .A2(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G190gat), .B(G218gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G134gat), .B(G162gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT36), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n460_));
  NAND2_X1  g259(.A1(G232gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G43gat), .B(G50gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(KEYINPUT15), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT15), .B1(new_n468_), .B2(new_n470_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT64), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n475_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT9), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT9), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G85gat), .A3(G92gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n486_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n481_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n490_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI211_X1 g299(.A(KEYINPUT8), .B(new_n496_), .C1(new_n500_), .C2(new_n486_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n503_));
  INV_X1    g302(.A(G99gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n475_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n484_), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n497_), .B(new_n505_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n496_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n502_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n495_), .B1(new_n501_), .B2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n474_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT68), .B1(new_n462_), .B2(new_n463_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n468_), .A2(new_n470_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n464_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n474_), .A2(new_n511_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n464_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n483_), .A2(new_n485_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n505_), .A2(new_n497_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n509_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT8), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n502_), .A3(new_n509_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n514_), .A3(new_n495_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n518_), .A2(new_n519_), .A3(new_n526_), .A4(new_n513_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n459_), .B1(new_n517_), .B2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n458_), .A2(KEYINPUT36), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n517_), .A2(new_n527_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n455_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G71gat), .B(G78gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(KEYINPUT11), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(G57gat), .ZN(new_n544_));
  INV_X1    g343(.A(G57gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G64gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n546_), .A3(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n541_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n511_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n495_), .B(new_n550_), .C1(new_n501_), .C2(new_n510_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(KEYINPUT65), .A3(new_n553_), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n511_), .A2(KEYINPUT65), .A3(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(G230gat), .ZN(new_n556_));
  INV_X1    g355(.A(G233gat), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(KEYINPUT12), .A3(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n511_), .A2(new_n561_), .A3(new_n551_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n538_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n558_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n553_), .A2(KEYINPUT12), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n550_), .B1(new_n525_), .B2(new_n495_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n562_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n537_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT13), .B1(new_n564_), .B2(new_n572_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT77), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n514_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n468_), .A2(KEYINPUT76), .A3(new_n470_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(KEYINPUT71), .A2(G15gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(KEYINPUT71), .A2(G15gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(G22gat), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(G22gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n588_), .B1(new_n589_), .B2(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT14), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT72), .B(G1gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n593_), .B2(G8gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT73), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(KEYINPUT72), .A2(G1gat), .ZN(new_n596_));
  NOR2_X1   g395(.A1(KEYINPUT72), .A2(G1gat), .ZN(new_n597_));
  OAI21_X1  g396(.A(G8gat), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT14), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n587_), .A4(new_n590_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G1gat), .B(G8gat), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n595_), .B2(new_n601_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n583_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n601_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n602_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n474_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n605_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n582_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT76), .B1(new_n468_), .B2(new_n470_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n611_), .B1(new_n605_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n579_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n611_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n603_), .A2(new_n583_), .A3(new_n604_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n615_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n579_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n605_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n575_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G127gat), .B(G155gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT16), .ZN(new_n629_));
  XOR2_X1   g428(.A(G183gat), .B(G211gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n550_), .B(KEYINPUT74), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n608_), .A2(new_n609_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(G231gat), .B(G233gat), .C1(new_n603_), .C2(new_n604_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n608_), .A2(new_n609_), .A3(new_n636_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n634_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT17), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n633_), .B1(new_n643_), .B2(new_n631_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT75), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n642_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n645_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n633_), .C1(new_n643_), .C2(new_n631_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n627_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n533_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n389_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G1gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n575_), .A2(KEYINPUT66), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n517_), .A2(new_n529_), .A3(new_n527_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT69), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT69), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n517_), .A2(new_n658_), .A3(new_n529_), .A4(new_n527_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n517_), .A2(new_n527_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n459_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n659_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT37), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT37), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT70), .B1(new_n531_), .B2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(new_n665_), .A3(new_n656_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT70), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT66), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n644_), .B(new_n648_), .ZN(new_n673_));
  AND4_X1   g472(.A1(new_n655_), .A2(new_n670_), .A3(new_n672_), .A4(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n399_), .A2(new_n422_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n427_), .A2(new_n428_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n452_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n453_), .A2(new_n454_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n674_), .B(new_n626_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT94), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n455_), .A2(KEYINPUT94), .A3(new_n626_), .A4(new_n674_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n388_), .A2(new_n593_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(KEYINPUT38), .A3(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n682_), .A3(new_n684_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n654_), .A2(new_n685_), .A3(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT95), .Z(G1324gat));
  NOR2_X1   g489(.A1(new_n427_), .A2(G8gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n681_), .A2(new_n682_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n681_), .A2(KEYINPUT96), .A3(new_n682_), .A4(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT98), .ZN(new_n697_));
  INV_X1    g496(.A(new_n427_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n455_), .A2(new_n698_), .A3(new_n532_), .A4(new_n651_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G8gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT39), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT39), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n702_), .A3(G8gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n697_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n697_), .B1(new_n696_), .B2(new_n704_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n706_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n696_), .A2(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT98), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n712_), .B2(new_n705_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1325gat));
  AOI21_X1  g513(.A(new_n438_), .B1(new_n652_), .B2(new_n452_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT41), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n683_), .A2(new_n438_), .A3(new_n452_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(KEYINPUT99), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(KEYINPUT99), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .ZN(G1326gat));
  INV_X1    g519(.A(new_n422_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n588_), .B1(new_n652_), .B2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT42), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n683_), .A2(new_n588_), .A3(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1327gat));
  OR2_X1    g524(.A1(new_n573_), .A2(new_n574_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT102), .B1(new_n673_), .B2(new_n532_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n650_), .A2(new_n728_), .A3(new_n531_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n455_), .A2(new_n730_), .A3(new_n626_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n731_), .A2(G29gat), .A3(new_n388_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n531_), .A2(KEYINPUT70), .A3(new_n665_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n667_), .A2(new_n668_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n733_), .A2(new_n734_), .B1(KEYINPUT37), .B2(new_n663_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n455_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT43), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n455_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n627_), .A2(new_n673_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(KEYINPUT44), .A3(new_n741_), .ZN(new_n742_));
  AOI211_X1 g541(.A(new_n673_), .B(new_n627_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n389_), .B(new_n742_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n745_), .A2(KEYINPUT101), .A3(G29gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT101), .B1(new_n745_), .B2(G29gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n732_), .B1(new_n746_), .B2(new_n747_), .ZN(G1328gat));
  NOR2_X1   g547(.A1(new_n427_), .A2(G36gat), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n455_), .A2(new_n730_), .A3(new_n626_), .A4(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n750_), .B(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(KEYINPUT46), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n698_), .B(new_n742_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G36gat), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n754_), .A2(KEYINPUT46), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1329gat));
  INV_X1    g558(.A(new_n452_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n435_), .B1(new_n731_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n452_), .A2(G43gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g564(.A1(new_n721_), .A2(G50gat), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n731_), .A2(new_n422_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n762_), .A2(new_n766_), .B1(G50gat), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(G1331gat));
  NOR3_X1   g569(.A1(new_n612_), .A2(new_n617_), .A3(new_n579_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n623_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n455_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT106), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n726_), .A2(new_n775_), .A3(new_n673_), .A4(new_n670_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n545_), .A3(new_n389_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n655_), .A2(new_n672_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n647_), .A2(new_n773_), .A3(new_n649_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n533_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n389_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n545_), .B2(new_n782_), .ZN(G1332gat));
  AOI21_X1  g582(.A(new_n543_), .B1(new_n781_), .B2(new_n698_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT48), .Z(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n543_), .A3(new_n698_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1333gat));
  INV_X1    g586(.A(G71gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n781_), .B2(new_n452_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT49), .Z(new_n790_));
  NAND3_X1  g589(.A1(new_n776_), .A2(new_n788_), .A3(new_n452_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1334gat));
  INV_X1    g591(.A(G78gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n781_), .B2(new_n721_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT50), .Z(new_n795_));
  NAND3_X1  g594(.A1(new_n776_), .A2(new_n793_), .A3(new_n721_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1335gat));
  NOR3_X1   g596(.A1(new_n673_), .A2(new_n626_), .A3(new_n575_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n740_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n389_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G85gat), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n727_), .A2(new_n729_), .B1(new_n655_), .B2(new_n672_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n775_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n389_), .A2(new_n487_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(G1336gat));
  OAI21_X1  g604(.A(new_n488_), .B1(new_n803_), .B2(new_n427_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n807_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n427_), .A2(new_n488_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n808_), .A2(new_n809_), .B1(new_n799_), .B2(new_n810_), .ZN(G1337gat));
  NAND2_X1  g610(.A1(new_n799_), .A2(new_n452_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G99gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n452_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n803_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g616(.A(new_n739_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n738_), .B1(new_n455_), .B2(new_n735_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n721_), .B(new_n798_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G106gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G106gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n721_), .A2(new_n475_), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n822_), .A2(new_n823_), .B1(new_n803_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR4_X1   g625(.A1(new_n735_), .A2(new_n779_), .A3(new_n726_), .A4(KEYINPUT54), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n735_), .A2(new_n726_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n780_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n611_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n605_), .A2(new_n610_), .A3(new_n619_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n578_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n578_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n835_), .A2(new_n836_), .B1(new_n564_), .B2(new_n572_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT55), .B1(new_n568_), .B2(new_n569_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n558_), .A2(KEYINPUT109), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n563_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n537_), .B1(new_n844_), .B2(new_n840_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n845_), .A3(KEYINPUT56), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT111), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  INV_X1    g647(.A(new_n842_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n844_), .B1(new_n570_), .B2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT55), .B(new_n840_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n538_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT110), .B(new_n848_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT111), .B1(new_n848_), .B2(KEYINPUT110), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n843_), .A2(new_n845_), .A3(new_n854_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n847_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n559_), .A2(new_n563_), .A3(new_n538_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT108), .B1(new_n773_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT108), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n572_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n838_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n862_), .B2(new_n532_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n848_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n846_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n857_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n865_), .A2(KEYINPUT58), .A3(new_n866_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n735_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT113), .B1(new_n863_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n532_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875_));
  INV_X1    g674(.A(new_n860_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n859_), .B1(new_n626_), .B2(new_n572_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n847_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n837_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n875_), .B1(new_n880_), .B2(new_n531_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n871_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n873_), .A2(new_n874_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n831_), .B1(new_n884_), .B2(new_n650_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n760_), .A2(new_n453_), .A3(new_n388_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT112), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(KEYINPUT112), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT114), .B1(new_n885_), .B2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n874_), .A2(new_n881_), .A3(new_n871_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n831_), .B1(new_n892_), .B2(new_n650_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n886_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT59), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n896_));
  INV_X1    g695(.A(new_n890_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n880_), .A2(new_n875_), .A3(new_n531_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n881_), .A2(new_n871_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(KEYINPUT113), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n673_), .B1(new_n900_), .B2(new_n883_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n896_), .B(new_n897_), .C1(new_n901_), .C2(new_n831_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n773_), .A2(new_n313_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n891_), .A2(new_n895_), .A3(new_n902_), .A4(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n893_), .A2(new_n894_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n313_), .B1(new_n906_), .B2(new_n773_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT115), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(new_n910_), .A3(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1340gat));
  XOR2_X1   g711(.A(KEYINPUT116), .B(G120gat), .Z(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n905_), .B(new_n914_), .C1(KEYINPUT60), .C2(new_n913_), .ZN(new_n915_));
  AND4_X1   g714(.A1(new_n778_), .A2(new_n891_), .A3(new_n895_), .A4(new_n902_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n913_), .ZN(G1341gat));
  NAND3_X1  g716(.A1(new_n905_), .A2(new_n308_), .A3(new_n673_), .ZN(new_n918_));
  AND4_X1   g717(.A1(new_n673_), .A2(new_n891_), .A3(new_n895_), .A4(new_n902_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n308_), .ZN(G1342gat));
  NAND3_X1  g719(.A1(new_n905_), .A2(new_n306_), .A3(new_n531_), .ZN(new_n921_));
  AND4_X1   g720(.A1(new_n735_), .A2(new_n891_), .A3(new_n895_), .A4(new_n902_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n306_), .ZN(G1343gat));
  NOR2_X1   g722(.A1(new_n452_), .A2(new_n422_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(new_n389_), .A3(new_n427_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n893_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n626_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n778_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT117), .B(G148gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1345gat));
  NAND2_X1  g730(.A1(new_n926_), .A2(new_n673_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n933_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1346gat));
  INV_X1    g739(.A(new_n926_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n670_), .ZN(new_n942_));
  INV_X1    g741(.A(G162gat), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n531_), .A2(new_n943_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n941_), .A2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT120), .B1(new_n944_), .B2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n948_));
  OAI221_X1 g747(.A(new_n948_), .B1(new_n941_), .B2(new_n945_), .C1(new_n942_), .C2(new_n943_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n454_), .A2(new_n427_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n422_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n626_), .B(new_n953_), .C1(new_n901_), .C2(new_n831_), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT122), .B1(new_n954_), .B2(G169gat), .ZN(new_n955_));
  XOR2_X1   g754(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n956_));
  OAI21_X1  g755(.A(KEYINPUT123), .B1(new_n885_), .B2(new_n952_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n958_), .B(new_n953_), .C1(new_n901_), .C2(new_n831_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n626_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(KEYINPUT124), .ZN(new_n962_));
  AOI22_X1  g761(.A1(new_n955_), .A2(new_n956_), .B1(new_n960_), .B2(new_n962_), .ZN(new_n963_));
  OR2_X1    g762(.A1(new_n955_), .A2(new_n956_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n954_), .A2(G169gat), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n963_), .B1(new_n964_), .B2(new_n967_), .ZN(G1348gat));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n892_), .A2(new_n650_), .ZN(new_n970_));
  OAI211_X1 g769(.A(new_n969_), .B(new_n422_), .C1(new_n970_), .C2(new_n831_), .ZN(new_n971_));
  OAI21_X1  g770(.A(KEYINPUT125), .B1(new_n893_), .B2(new_n721_), .ZN(new_n972_));
  NAND4_X1  g771(.A1(new_n971_), .A2(new_n972_), .A3(new_n778_), .A4(new_n951_), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n973_), .A2(G176gat), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n575_), .A2(G176gat), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n976_), .B1(new_n957_), .B2(new_n959_), .ZN(new_n977_));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n974_), .B2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n973_), .A2(G176gat), .ZN(new_n980_));
  AND2_X1   g779(.A1(new_n957_), .A2(new_n959_), .ZN(new_n981_));
  OAI211_X1 g780(.A(new_n979_), .B(new_n980_), .C1(new_n981_), .C2(new_n976_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n978_), .A2(new_n982_), .ZN(G1349gat));
  NAND3_X1  g782(.A1(new_n971_), .A2(new_n972_), .A3(new_n951_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(new_n650_), .ZN(new_n985_));
  AOI21_X1  g784(.A(G183gat), .B1(new_n985_), .B2(KEYINPUT127), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n987_), .B1(new_n984_), .B2(new_n650_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n650_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n989_));
  AOI22_X1  g788(.A1(new_n986_), .A2(new_n988_), .B1(new_n960_), .B2(new_n989_), .ZN(G1350gat));
  OAI21_X1  g789(.A(G190gat), .B1(new_n981_), .B2(new_n670_), .ZN(new_n991_));
  NAND3_X1  g790(.A1(new_n531_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n992_));
  OAI21_X1  g791(.A(new_n991_), .B1(new_n981_), .B2(new_n992_), .ZN(G1351gat));
  NAND3_X1  g792(.A1(new_n924_), .A2(new_n388_), .A3(new_n698_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(new_n893_), .A2(new_n994_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n995_), .A2(new_n626_), .ZN(new_n996_));
  XNOR2_X1  g795(.A(new_n996_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g796(.A1(new_n995_), .A2(new_n778_), .ZN(new_n998_));
  XNOR2_X1  g797(.A(new_n998_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g798(.A1(new_n995_), .A2(new_n673_), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1001_));
  AND2_X1   g800(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1002_));
  NOR3_X1   g801(.A1(new_n1000_), .A2(new_n1001_), .A3(new_n1002_), .ZN(new_n1003_));
  AOI21_X1  g802(.A(new_n1003_), .B1(new_n1000_), .B2(new_n1001_), .ZN(G1354gat));
  NAND3_X1  g803(.A1(new_n995_), .A2(new_n255_), .A3(new_n531_), .ZN(new_n1005_));
  NOR3_X1   g804(.A1(new_n893_), .A2(new_n670_), .A3(new_n994_), .ZN(new_n1006_));
  OAI21_X1  g805(.A(new_n1005_), .B1(new_n1006_), .B2(new_n255_), .ZN(G1355gat));
endmodule


