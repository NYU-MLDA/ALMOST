//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT0), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G57gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n204_), .A2(new_n205_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n205_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(G85gat), .A3(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G225gat), .A2(G233gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G127gat), .B(G134gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  AND3_X1   g015(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n226_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n229_), .B(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n216_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n213_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n214_), .B(new_n215_), .Z(new_n244_));
  INV_X1    g043(.A(new_n232_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n222_), .A2(new_n224_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n226_), .B1(new_n246_), .B2(KEYINPUT1), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n247_), .B2(new_n225_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n227_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n231_), .B(KEYINPUT3), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n229_), .B(KEYINPUT2), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n244_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT100), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n233_), .A2(new_n216_), .A3(new_n239_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n233_), .A2(new_n239_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT100), .A3(new_n244_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n243_), .B1(new_n259_), .B2(KEYINPUT4), .ZN(new_n260_));
  INV_X1    g059(.A(new_n213_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n212_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n213_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n208_), .A2(new_n211_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n241_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n264_), .B(new_n265_), .C1(new_n266_), .C2(new_n243_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270_));
  INV_X1    g069(.A(G204gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(G197gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(G197gat), .ZN(new_n273_));
  INV_X1    g072(.A(G197gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n272_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277_));
  INV_X1    g076(.A(G211gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(G218gat), .ZN(new_n279_));
  INV_X1    g078(.A(G218gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(G211gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT91), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(G211gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(G218gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n276_), .A2(new_n277_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G197gat), .B(G204gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT89), .B1(new_n288_), .B2(new_n277_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n274_), .A2(G204gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n273_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT21), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n286_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n285_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n272_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n298_), .A2(KEYINPUT21), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n287_), .A2(new_n294_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G233gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(G228gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(G228gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n300_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n257_), .A2(KEYINPUT29), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT92), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT92), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(new_n311_), .A3(new_n308_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT93), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n257_), .A2(KEYINPUT93), .A3(KEYINPUT29), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n282_), .A2(new_n298_), .A3(KEYINPUT21), .A4(new_n286_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n292_), .B1(new_n291_), .B2(KEYINPUT21), .ZN(new_n317_));
  AOI211_X1 g116(.A(KEYINPUT89), .B(new_n277_), .C1(new_n273_), .C2(new_n290_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n295_), .A2(new_n296_), .B1(new_n298_), .B2(KEYINPUT21), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n315_), .A3(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n310_), .A2(new_n312_), .B1(new_n322_), .B2(new_n306_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT94), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n257_), .A2(KEYINPUT29), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT87), .ZN(new_n328_));
  XOR2_X1   g127(.A(G22gat), .B(G50gat), .Z(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT28), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n310_), .A2(new_n312_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n322_), .A2(new_n306_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(new_n324_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n323_), .A2(new_n325_), .ZN(new_n336_));
  OAI22_X1  g135(.A1(new_n326_), .A2(new_n331_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n329_), .B(KEYINPUT28), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n328_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n324_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n323_), .A2(new_n325_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT94), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n344_));
  INV_X1    g143(.A(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT24), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT23), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G183gat), .A3(G190gat), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT79), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(G190gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT26), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n362_), .B2(new_n356_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G183gat), .ZN(new_n365_));
  INV_X1    g164(.A(G183gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT25), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n367_), .A3(KEYINPUT76), .ZN(new_n368_));
  OR3_X1    g167(.A1(new_n366_), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT24), .ZN(new_n372_));
  INV_X1    g171(.A(new_n348_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n351_), .A2(new_n353_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n347_), .A2(KEYINPUT24), .A3(new_n348_), .A4(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n355_), .A2(new_n371_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT81), .B(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n346_), .B1(new_n383_), .B2(KEYINPUT80), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n382_), .B(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n353_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n351_), .A2(new_n353_), .A3(new_n387_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n381_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n321_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G169gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n346_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n379_), .B(KEYINPUT97), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n395_), .B(new_n396_), .C1(new_n354_), .C2(new_n386_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n375_), .A2(new_n388_), .A3(new_n380_), .A4(new_n389_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n359_), .A2(new_n361_), .A3(KEYINPUT96), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT96), .B1(new_n359_), .B2(new_n361_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n365_), .A2(new_n367_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT99), .B1(new_n321_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT99), .ZN(new_n405_));
  INV_X1    g204(.A(new_n390_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT96), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n362_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n359_), .A2(new_n361_), .A3(KEYINPUT96), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n408_), .A2(new_n365_), .A3(new_n367_), .A4(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n406_), .A2(new_n410_), .A3(new_n375_), .A4(new_n380_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n300_), .A2(new_n405_), .A3(new_n411_), .A4(new_n397_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n393_), .A2(new_n404_), .A3(new_n412_), .A4(KEYINPUT20), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT95), .Z(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT19), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n381_), .A2(new_n391_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n300_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n416_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT98), .B1(new_n321_), .B2(new_n403_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n321_), .A2(new_n403_), .A3(KEYINPUT98), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT18), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G64gat), .ZN(new_n428_));
  INV_X1    g227(.A(G92gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n417_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(KEYINPUT27), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n404_), .A2(new_n412_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n418_), .B1(new_n392_), .B2(new_n321_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n421_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n321_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n321_), .A2(new_n403_), .A3(KEYINPUT98), .ZN(new_n440_));
  NOR4_X1   g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n422_), .A4(new_n416_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n430_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n442_));
  NOR4_X1   g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n422_), .A4(new_n421_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n300_), .A2(new_n397_), .A3(new_n411_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n416_), .B1(new_n437_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n431_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n442_), .A2(new_n446_), .A3(KEYINPUT27), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n343_), .A2(new_n435_), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G15gat), .B(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT84), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT83), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n450_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n419_), .A2(KEYINPUT30), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n392_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT31), .ZN(new_n461_));
  INV_X1    g260(.A(new_n459_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(new_n457_), .A3(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n454_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n463_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT31), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n453_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n466_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n216_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n466_), .A2(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT85), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n466_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n244_), .A3(new_n477_), .ZN(new_n478_));
  AND4_X1   g277(.A1(new_n269_), .A2(new_n448_), .A3(new_n474_), .A4(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n255_), .A2(new_n254_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(new_n240_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n258_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT4), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n262_), .B1(new_n484_), .B2(new_n242_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT33), .B1(new_n485_), .B2(new_n265_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487_));
  NOR4_X1   g286(.A1(new_n260_), .A2(new_n487_), .A3(new_n212_), .A4(new_n262_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n261_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT101), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n212_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n213_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT101), .B1(new_n493_), .B2(new_n265_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n261_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n484_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n489_), .A2(new_n434_), .A3(KEYINPUT102), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT102), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n417_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n442_), .A2(new_n500_), .A3(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n267_), .A2(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n484_), .A2(new_n242_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n503_), .A2(KEYINPUT33), .A3(new_n264_), .A4(new_n265_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n499_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n443_), .A2(new_n445_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n268_), .B(new_n508_), .C1(new_n509_), .C2(new_n507_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n498_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n343_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n511_), .A2(KEYINPUT103), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT103), .B1(new_n511_), .B2(new_n512_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n435_), .A2(new_n447_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n269_), .A3(new_n343_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n513_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n474_), .A2(new_n478_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n480_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(G22gat), .ZN(new_n522_));
  INV_X1    g321(.A(G15gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT73), .B(G8gat), .Z(new_n525_));
  INV_X1    g324(.A(G1gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G1gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G8gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(G8gat), .A3(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G29gat), .B(G36gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n538_), .B(KEYINPUT15), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT75), .B1(new_n535_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n542_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n539_), .B(new_n540_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n535_), .B(new_n538_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n540_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G169gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n274_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n546_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT10), .B(G99gat), .Z(new_n561_));
  INV_X1    g360(.A(G106gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G85gat), .B(G92gat), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT9), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n207_), .A2(new_n429_), .A3(KEYINPUT9), .ZN(new_n566_));
  AND3_X1   g365(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n563_), .A2(new_n565_), .A3(new_n566_), .A4(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT64), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT65), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT7), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT65), .ZN(new_n579_));
  NOR2_X1   g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n575_), .A2(new_n569_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n564_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT8), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT8), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n564_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT66), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n575_), .A2(KEYINPUT66), .A3(new_n581_), .A4(new_n569_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n584_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  AOI211_X1 g391(.A(KEYINPUT67), .B(new_n586_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n570_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT68), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT11), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n598_), .B2(new_n597_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(KEYINPUT11), .A3(new_n595_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n594_), .A2(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n603_), .B(new_n570_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(KEYINPUT12), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n594_), .A2(new_n608_), .A3(new_n604_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n560_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n559_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n271_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT5), .B(G176gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n610_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT70), .B1(new_n617_), .B2(KEYINPUT69), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n607_), .A2(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n559_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n611_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n615_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT69), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT70), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n615_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n618_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n618_), .B2(new_n625_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n558_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n618_), .A2(new_n625_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n618_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(KEYINPUT13), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n594_), .A2(new_n541_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT34), .ZN(new_n639_));
  INV_X1    g438(.A(new_n538_), .ZN(new_n640_));
  OAI221_X1 g439(.A(new_n637_), .B1(KEYINPUT35), .B2(new_n639_), .C1(new_n640_), .C2(new_n594_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(KEYINPUT35), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT71), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n641_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G190gat), .B(G218gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G134gat), .B(G162gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT36), .Z(new_n648_));
  AND2_X1   g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(KEYINPUT36), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n644_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n636_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n644_), .A2(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n644_), .A2(new_n648_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(KEYINPUT37), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n535_), .B(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(new_n603_), .ZN(new_n660_));
  XOR2_X1   g459(.A(G183gat), .B(G211gat), .Z(new_n661_));
  XNOR2_X1  g460(.A(G127gat), .B(G155gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT17), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n660_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n660_), .A2(KEYINPUT17), .A3(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n657_), .A2(new_n669_), .ZN(new_n670_));
  AND4_X1   g469(.A1(new_n521_), .A2(new_n557_), .A3(new_n635_), .A4(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n526_), .A3(new_n268_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT104), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT38), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n654_), .A2(new_n655_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n521_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n557_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n635_), .ZN(new_n678_));
  NOR4_X1   g477(.A1(new_n676_), .A2(new_n669_), .A3(new_n677_), .A4(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n526_), .B1(new_n679_), .B2(new_n268_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT105), .Z(new_n681_));
  NAND2_X1  g480(.A1(new_n674_), .A2(new_n681_), .ZN(G1324gat));
  INV_X1    g481(.A(new_n515_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n671_), .A2(new_n683_), .A3(new_n525_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n679_), .A2(new_n683_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G8gat), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  NAND3_X1  g490(.A1(new_n671_), .A2(new_n523_), .A3(new_n520_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT106), .Z(new_n693_));
  AOI21_X1  g492(.A(new_n523_), .B1(new_n679_), .B2(new_n520_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  INV_X1    g497(.A(G22gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n679_), .B2(new_n343_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n671_), .A2(new_n699_), .A3(new_n343_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(new_n675_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n521_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n635_), .A2(new_n669_), .A3(new_n557_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n268_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n657_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n521_), .A2(new_n657_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n511_), .A2(new_n512_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n511_), .A2(KEYINPUT103), .A3(new_n512_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n516_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n479_), .B1(new_n719_), .B2(new_n519_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n657_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n712_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n707_), .B1(new_n714_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT44), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(G29gat), .A3(new_n268_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n714_), .A2(new_n722_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n707_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT109), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n713_), .B1(new_n521_), .B2(new_n657_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n720_), .A2(new_n721_), .A3(new_n712_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n732_), .B(new_n727_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n729_), .A2(new_n731_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n709_), .B1(new_n725_), .B2(new_n736_), .ZN(G1328gat));
  AOI21_X1  g536(.A(new_n515_), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n731_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n723_), .A2(new_n732_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT111), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n738_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(G36gat), .A3(new_n744_), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n706_), .A2(new_n707_), .A3(G36gat), .A4(new_n515_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT45), .Z(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(KEYINPUT46), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1329gat));
  NAND3_X1  g551(.A1(new_n736_), .A2(new_n520_), .A3(new_n724_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n519_), .A2(G43gat), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n753_), .A2(G43gat), .B1(new_n708_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1330gat));
  AOI21_X1  g556(.A(G50gat), .B1(new_n708_), .B2(new_n343_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n736_), .A2(new_n724_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n343_), .A2(G50gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n678_), .A2(new_n670_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT113), .Z(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n720_), .A3(new_n557_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n205_), .A3(new_n268_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n678_), .A2(new_n677_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n676_), .A2(new_n766_), .A3(new_n669_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G57gat), .B1(new_n768_), .B2(new_n269_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(G1332gat));
  INV_X1    g569(.A(G64gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n767_), .B2(new_n683_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT48), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n683_), .A2(new_n771_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT114), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n764_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n767_), .B2(new_n520_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT49), .Z(new_n780_));
  NAND3_X1  g579(.A1(new_n764_), .A2(new_n778_), .A3(new_n520_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1334gat));
  INV_X1    g581(.A(G78gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n767_), .B2(new_n343_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT50), .Z(new_n785_));
  NAND3_X1  g584(.A1(new_n764_), .A2(new_n783_), .A3(new_n343_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1335gat));
  NAND3_X1  g586(.A1(new_n678_), .A2(new_n669_), .A3(new_n677_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n790_), .A2(new_n791_), .B1(new_n714_), .B2(new_n722_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793_), .B2(new_n269_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n706_), .A2(new_n788_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n207_), .A3(new_n268_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n793_), .B2(new_n515_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n429_), .A3(new_n683_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n793_), .B2(new_n519_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n795_), .A2(new_n520_), .A3(new_n561_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(KEYINPUT116), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n803_), .B(new_n805_), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n795_), .A2(new_n562_), .A3(new_n343_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n792_), .A2(new_n343_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(G106gat), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT52), .B(new_n562_), .C1(new_n792_), .C2(new_n343_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g612(.A1(new_n657_), .A2(new_n669_), .A3(new_n557_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n635_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n814_), .B2(new_n635_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n547_), .A2(new_n540_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n554_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n539_), .A2(new_n548_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n545_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n543_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT120), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n539_), .B(new_n548_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n554_), .A4(new_n820_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(new_n556_), .A3(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n627_), .A2(new_n628_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n620_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n619_), .A2(KEYINPUT118), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n607_), .A2(new_n835_), .A3(new_n609_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n560_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT55), .B1(new_n610_), .B2(KEYINPUT117), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT119), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n839_), .B2(new_n616_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n839_), .A2(new_n844_), .A3(KEYINPUT56), .A4(new_n616_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n677_), .A2(new_n617_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n830_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n819_), .B1(new_n848_), .B2(new_n705_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n847_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n839_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n842_), .B1(new_n851_), .B2(new_n844_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n841_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT57), .B(new_n675_), .C1(new_n853_), .C2(new_n830_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n851_), .A2(new_n842_), .A3(KEYINPUT121), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n829_), .A2(new_n617_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n839_), .A2(KEYINPUT121), .A3(KEYINPUT56), .A4(new_n616_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n843_), .A2(new_n861_), .A3(new_n840_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n862_), .A2(KEYINPUT58), .A3(new_n858_), .A4(new_n857_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n863_), .A3(new_n657_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n849_), .A2(new_n854_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n818_), .B1(new_n865_), .B2(new_n669_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n519_), .A2(new_n269_), .A3(new_n343_), .A4(new_n683_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT122), .Z(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n557_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  INV_X1    g672(.A(new_n669_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n675_), .B1(new_n853_), .B2(new_n830_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n840_), .A2(new_n861_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n859_), .B1(new_n876_), .B2(new_n843_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n721_), .B1(new_n877_), .B2(KEYINPUT58), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n875_), .A2(new_n819_), .B1(new_n878_), .B2(new_n860_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n874_), .B1(new_n879_), .B2(new_n854_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n873_), .B(new_n868_), .C1(new_n880_), .C2(new_n818_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n866_), .B2(new_n869_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n557_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n872_), .B1(new_n883_), .B2(new_n871_), .ZN(G1340gat));
  AND3_X1   g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n678_), .ZN(new_n885_));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n870_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n635_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(KEYINPUT60), .B2(new_n886_), .ZN(new_n889_));
  OAI22_X1  g688(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n889_), .ZN(G1341gat));
  NAND3_X1  g689(.A1(new_n881_), .A2(new_n882_), .A3(new_n874_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G127gat), .ZN(new_n892_));
  INV_X1    g691(.A(G127gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n870_), .A2(new_n893_), .A3(new_n874_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT123), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n897_), .A3(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1342gat));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n870_), .A2(new_n900_), .A3(new_n705_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n881_), .A2(new_n882_), .A3(new_n657_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n900_), .ZN(G1343gat));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  INV_X1    g703(.A(new_n866_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n683_), .A2(new_n512_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n519_), .A2(new_n906_), .A3(new_n268_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n866_), .A2(KEYINPUT124), .A3(new_n907_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n557_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g711(.A(new_n678_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g713(.A(new_n874_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1346gat));
  OR2_X1    g716(.A1(new_n909_), .A2(new_n910_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n657_), .A2(G162gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT125), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n705_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n921_));
  INV_X1    g720(.A(G162gat), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n918_), .A2(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1347gat));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n519_), .A2(new_n268_), .A3(new_n343_), .A4(new_n515_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n905_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n677_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n924_), .B1(new_n927_), .B2(new_n345_), .ZN(new_n928_));
  OAI211_X1 g727(.A(KEYINPUT62), .B(G169gat), .C1(new_n926_), .C2(new_n677_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n394_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(G1348gat));
  NOR2_X1   g730(.A1(new_n926_), .A2(new_n635_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n346_), .ZN(G1349gat));
  NOR2_X1   g732(.A1(new_n926_), .A2(new_n669_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(G183gat), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n401_), .B2(new_n934_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n926_), .B2(new_n721_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n705_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n926_), .B2(new_n938_), .ZN(G1351gat));
  NOR4_X1   g738(.A1(new_n520_), .A2(new_n268_), .A3(new_n512_), .A4(new_n515_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n905_), .A2(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n677_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n274_), .ZN(G1352gat));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n635_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT126), .B(G204gat), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1353gat));
  INV_X1    g745(.A(new_n941_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n874_), .B1(new_n948_), .B2(new_n278_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT127), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n947_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n948_), .A2(new_n278_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n941_), .B2(new_n721_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n705_), .A2(new_n280_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n941_), .B2(new_n955_), .ZN(G1355gat));
endmodule


