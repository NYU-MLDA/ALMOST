//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT76), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT36), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  AND2_X1   g013(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NOR4_X1   g018(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT64), .A4(G106gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n213_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G85gat), .B2(G92gat), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G85gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT66), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G92gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT9), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n223_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT67), .B1(new_n221_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n223_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n225_), .A2(new_n227_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(KEYINPUT9), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT10), .B(G99gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(new_n241_), .B2(G106gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n217_), .A2(new_n214_), .A3(new_n218_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n240_), .A2(new_n244_), .A3(new_n245_), .A4(new_n213_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  INV_X1    g046(.A(G99gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n218_), .A3(KEYINPUT69), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(G99gat), .B2(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT68), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n256_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n253_), .A2(new_n255_), .A3(new_n213_), .A4(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n224_), .A2(new_n229_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G85gat), .A2(G92gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n247_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n247_), .A3(new_n261_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n237_), .B(new_n246_), .C1(new_n262_), .C2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G29gat), .B(G36gat), .Z(new_n266_));
  XOR2_X1   g065(.A(G43gat), .B(G50gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT34), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n271_), .A2(KEYINPUT35), .ZN(new_n272_));
  INV_X1    g071(.A(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT15), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT15), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n268_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n265_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n269_), .A2(new_n272_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n269_), .A2(KEYINPUT75), .A3(new_n272_), .A4(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n269_), .A2(new_n278_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n271_), .A2(KEYINPUT35), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n272_), .A2(new_n284_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n281_), .A2(new_n282_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n206_), .A2(new_n207_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n208_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(KEYINPUT77), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(new_n282_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n285_), .ZN(new_n292_));
  AOI221_X4 g091(.A(KEYINPUT77), .B1(new_n208_), .B2(new_n287_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT78), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n202_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n288_), .B(new_n289_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(KEYINPUT78), .A3(KEYINPUT37), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT13), .ZN(new_n300_));
  INV_X1    g099(.A(new_n262_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n263_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G64gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n305_));
  XOR2_X1   g104(.A(G71gat), .B(G78gat), .Z(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n302_), .A2(new_n309_), .A3(new_n237_), .A4(new_n246_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G230gat), .A2(G233gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT70), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT12), .ZN(new_n313_));
  INV_X1    g112(.A(new_n309_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n265_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n265_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT70), .B1(new_n310_), .B2(new_n311_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT71), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n265_), .A2(new_n314_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n310_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G230gat), .A3(G233gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(KEYINPUT12), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n265_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n310_), .A2(new_n311_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n325_), .A2(new_n328_), .A3(new_n329_), .A4(new_n312_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n319_), .A2(new_n322_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G176gat), .B(G204gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT73), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n319_), .A2(new_n322_), .A3(new_n330_), .A4(new_n337_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT74), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT74), .B1(new_n339_), .B2(new_n340_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n300_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n340_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(KEYINPUT13), .A3(new_n341_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G231gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n309_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT79), .B(G1gat), .ZN(new_n352_));
  INV_X1    g151(.A(G8gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT14), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G15gat), .B(G22gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G8gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n351_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT80), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G155gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT16), .ZN(new_n365_));
  XOR2_X1   g164(.A(G183gat), .B(G211gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT17), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n363_), .B(new_n369_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n362_), .A2(KEYINPUT17), .A3(new_n368_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n299_), .A2(new_n349_), .A3(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT81), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n273_), .B1(new_n360_), .B2(new_n359_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n274_), .A2(new_n360_), .A3(new_n359_), .A4(new_n276_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G229gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT82), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n361_), .B(new_n268_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G229gat), .A3(G233gat), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT83), .A4(new_n380_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G141gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G169gat), .B(G197gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .A4(new_n390_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT84), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n387_), .A2(new_n395_), .A3(new_n391_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT88), .B(G176gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT22), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(G169gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n400_), .B(new_n403_), .C1(new_n404_), .C2(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT23), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n399_), .B(new_n405_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n399_), .A2(KEYINPUT24), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  MUX2_X1   g215(.A(new_n415_), .B(KEYINPUT24), .S(new_n416_), .Z(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT25), .B(G183gat), .ZN(new_n418_));
  INV_X1    g217(.A(G190gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT26), .B1(new_n419_), .B2(KEYINPUT85), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(KEYINPUT26), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n418_), .B(new_n420_), .C1(new_n421_), .C2(KEYINPUT85), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n410_), .B1(G183gat), .B2(G190gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G127gat), .B(G134gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT91), .ZN(new_n434_));
  XOR2_X1   g233(.A(G113gat), .B(G120gat), .Z(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n434_), .B(new_n435_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n432_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n431_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n429_), .A2(new_n430_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(G43gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G15gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n447_), .A2(KEYINPUT31), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(KEYINPUT31), .ZN(new_n449_));
  OR3_X1    g248(.A1(new_n440_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n440_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G211gat), .B(G218gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT21), .ZN(new_n458_));
  INV_X1    g257(.A(G204gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G197gat), .ZN(new_n460_));
  INV_X1    g259(.A(G197gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G204gat), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n458_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(KEYINPUT94), .A3(G197gat), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n458_), .A4(new_n462_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n468_), .A2(KEYINPUT95), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(KEYINPUT95), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n467_), .A3(new_n462_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n457_), .A2(KEYINPUT21), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G141gat), .A2(G148gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT3), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G141gat), .A2(G148gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT2), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(KEYINPUT1), .B2(new_n481_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(KEYINPUT1), .B2(new_n481_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n476_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n487_), .A2(new_n478_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n480_), .A2(new_n484_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n474_), .B1(new_n475_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(KEYINPUT93), .A2(G233gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT93), .A2(G233gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(G228gat), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(new_n495_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n454_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n454_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n475_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G22gat), .B(G50gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT28), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n502_), .B(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n498_), .B2(KEYINPUT97), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n499_), .A2(KEYINPUT97), .A3(new_n500_), .A4(new_n505_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G225gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n434_), .A2(new_n435_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n434_), .A2(new_n435_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n432_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n489_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n436_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n489_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT100), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n437_), .A2(new_n522_), .A3(new_n489_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n438_), .A2(KEYINPUT99), .A3(new_n515_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n511_), .B(new_n519_), .C1(new_n528_), .C2(new_n518_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n521_), .A2(new_n523_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT99), .B1(new_n438_), .B2(new_n515_), .ZN(new_n531_));
  AND4_X1   g330(.A1(KEYINPUT99), .A2(new_n514_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n510_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G1gat), .B(G29gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G85gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(KEYINPUT33), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT102), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT102), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT33), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n540_), .B1(new_n528_), .B2(new_n511_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n519_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n533_), .B2(KEYINPUT4), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n550_), .B2(new_n511_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT103), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G8gat), .B(G36gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT18), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G64gat), .B(G92gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G226gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT19), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n471_), .A2(new_n414_), .A3(new_n473_), .A4(new_n426_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(KEYINPUT20), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n404_), .A2(new_n400_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n399_), .B(new_n564_), .C1(new_n425_), .C2(new_n413_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n418_), .ZN(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT26), .B(G190gat), .Z(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n568_), .A2(new_n411_), .A3(new_n409_), .A4(new_n417_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n474_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n561_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n570_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n474_), .A2(new_n427_), .ZN(new_n575_));
  AND4_X1   g374(.A1(KEYINPUT20), .A2(new_n574_), .A3(new_n575_), .A4(new_n561_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n558_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n579_));
  INV_X1    g378(.A(new_n474_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n573_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n561_), .A3(new_n575_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n571_), .A2(KEYINPUT20), .A3(new_n562_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n560_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n584_), .A3(new_n557_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n578_), .A3(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n582_), .A2(new_n584_), .A3(KEYINPUT98), .A4(new_n557_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT103), .B(new_n548_), .C1(new_n550_), .C2(new_n511_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n553_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n528_), .A2(new_n511_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n550_), .B2(new_n511_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n593_), .B2(new_n543_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n547_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n543_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n544_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n561_), .B1(new_n581_), .B2(new_n575_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n583_), .A2(new_n560_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n557_), .A2(KEYINPUT32), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n582_), .A2(new_n602_), .A3(new_n584_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n509_), .B1(new_n595_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n598_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n509_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n586_), .A2(new_n587_), .A3(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT27), .B(new_n585_), .C1(new_n601_), .C2(new_n557_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n452_), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n452_), .A2(new_n598_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n509_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n612_), .A2(KEYINPUT105), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n612_), .A2(KEYINPUT105), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n615_), .B(new_n616_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n398_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n374_), .A2(KEYINPUT81), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n375_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n598_), .A3(new_n352_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n297_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n349_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n397_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n373_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n607_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n624_), .A2(new_n625_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n633_), .A3(new_n634_), .ZN(G1324gat));
  NOR2_X1   g434(.A1(new_n617_), .A2(new_n618_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n623_), .A2(new_n353_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n638_), .B2(KEYINPUT106), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n631_), .B2(new_n636_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n640_), .A2(KEYINPUT106), .A3(new_n638_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(KEYINPUT106), .B2(new_n638_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n637_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT40), .B(new_n637_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1325gat));
  OAI21_X1  g446(.A(G15gat), .B1(new_n632_), .B2(new_n452_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT41), .Z(new_n649_));
  NOR3_X1   g448(.A1(new_n622_), .A2(G15gat), .A3(new_n452_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT107), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(G1326gat));
  OAI21_X1  g451(.A(G22gat), .B1(new_n632_), .B2(new_n616_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n616_), .A2(G22gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n622_), .B2(new_n655_), .ZN(G1327gat));
  NOR3_X1   g455(.A1(new_n349_), .A2(new_n372_), .A3(new_n294_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n620_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n598_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n299_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n296_), .A2(new_n298_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT108), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n299_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n452_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT33), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n545_), .B1(new_n544_), .B2(KEYINPUT33), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n594_), .A2(new_n588_), .A3(new_n589_), .A4(new_n553_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n605_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n616_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n608_), .A2(new_n612_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n619_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n666_), .B(new_n668_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n664_), .B1(new_n679_), .B2(KEYINPUT43), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n629_), .A2(new_n372_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n661_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n299_), .B(KEYINPUT108), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n614_), .A2(new_n619_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n662_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n681_), .C1(new_n686_), .C2(new_n664_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n683_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n598_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n660_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n636_), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n636_), .A2(KEYINPUT109), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n636_), .A2(KEYINPUT109), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n658_), .A2(G36gat), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT111), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n697_), .B(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n692_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n692_), .A2(KEYINPUT46), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND4_X1  g504(.A1(new_n683_), .A2(G43gat), .A3(new_n687_), .A4(new_n669_), .ZN(new_n706_));
  INV_X1    g505(.A(G43gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n658_), .B2(new_n452_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g509(.A(G50gat), .B1(new_n659_), .B2(new_n509_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n509_), .A2(G50gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n688_), .B2(new_n712_), .ZN(G1331gat));
  AOI211_X1 g512(.A(new_n397_), .B(new_n628_), .C1(new_n614_), .C2(new_n619_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n299_), .A2(new_n373_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n598_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n628_), .A2(new_n397_), .A3(new_n373_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n627_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n607_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n720_), .B2(new_n696_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n696_), .A2(G64gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT112), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n716_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1333gat));
  NOR2_X1   g527(.A1(new_n452_), .A2(G71gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n716_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n627_), .A2(new_n669_), .A3(new_n719_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G71gat), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT49), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT49), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT114), .Z(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n720_), .B2(new_n616_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT50), .ZN(new_n739_));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n716_), .A2(new_n740_), .A3(new_n509_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1335gat));
  NAND3_X1  g541(.A1(new_n349_), .A2(new_n398_), .A3(new_n373_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT116), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n680_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n598_), .A3(new_n228_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n294_), .A2(new_n372_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n714_), .A2(new_n598_), .A3(new_n747_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n748_), .A2(KEYINPUT115), .A3(new_n224_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT115), .B1(new_n748_), .B2(new_n224_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1336gat));
  NAND2_X1  g552(.A1(new_n714_), .A2(new_n747_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G92gat), .B1(new_n755_), .B2(new_n636_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n695_), .A2(new_n233_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n745_), .B2(new_n757_), .ZN(G1337gat));
  AOI21_X1  g557(.A(new_n248_), .B1(new_n745_), .B2(new_n669_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n754_), .A2(new_n452_), .A3(new_n241_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(KEYINPUT118), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n761_), .B(new_n764_), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n755_), .A2(new_n218_), .A3(new_n509_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n743_), .B(KEYINPUT116), .Z(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n509_), .C1(new_n686_), .C2(new_n664_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n766_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n766_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n390_), .B1(new_n384_), .B2(new_n380_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n377_), .A2(new_n378_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n380_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n393_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n347_), .B2(new_n341_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n397_), .A2(new_n340_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n319_), .A2(new_n785_), .A3(new_n330_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT119), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n319_), .A2(new_n788_), .A3(new_n330_), .A4(new_n785_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n310_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(G230gat), .A3(G233gat), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n325_), .A2(new_n328_), .A3(KEYINPUT55), .A4(new_n312_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n787_), .A2(new_n789_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n338_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n784_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n793_), .B1(new_n786_), .B2(KEYINPUT119), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n337_), .B1(new_n800_), .B2(new_n789_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n797_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n783_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n777_), .B1(new_n803_), .B2(new_n297_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n781_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n397_), .B(new_n340_), .C1(new_n801_), .C2(new_n797_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n796_), .A2(new_n798_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n294_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n801_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n340_), .A2(new_n781_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n801_), .B2(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n812_), .A3(KEYINPUT58), .A4(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n299_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n804_), .A2(new_n809_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n804_), .A2(new_n819_), .A3(new_n809_), .A4(KEYINPUT121), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n373_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n715_), .A2(new_n398_), .A3(new_n628_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT54), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n374_), .A2(new_n827_), .A3(new_n398_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n636_), .A2(new_n509_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n598_), .A3(new_n669_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n397_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n820_), .A2(new_n373_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n833_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n398_), .A2(new_n835_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n832_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n840_), .B(new_n841_), .C1(new_n842_), .C2(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT122), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n836_), .A2(new_n843_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n628_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n842_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n349_), .B(new_n840_), .C1(new_n842_), .C2(new_n839_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n853_), .B2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n842_), .B2(new_n372_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(KEYINPUT123), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(KEYINPUT123), .ZN(new_n857_));
  INV_X1    g656(.A(new_n840_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n842_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(KEYINPUT59), .B2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n372_), .A2(G127gat), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n856_), .A2(new_n857_), .B1(new_n860_), .B2(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n842_), .B2(new_n297_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT124), .B(G134gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n665_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n860_), .B2(new_n865_), .ZN(G1343gat));
  AOI21_X1  g665(.A(new_n669_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n695_), .A2(new_n607_), .A3(new_n616_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n398_), .ZN(new_n870_));
  INV_X1    g669(.A(G141gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n628_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT125), .B(G148gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  NOR2_X1   g674(.A1(new_n869_), .A2(new_n373_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n876_), .B(new_n878_), .ZN(G1346gat));
  AND2_X1   g678(.A1(new_n867_), .A2(new_n868_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G162gat), .B1(new_n880_), .B2(new_n297_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n684_), .A2(G162gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(new_n882_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n695_), .A2(new_n616_), .A3(new_n615_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n838_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n398_), .ZN(new_n887_));
  INV_X1    g686(.A(G169gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n404_), .ZN(new_n890_));
  OAI211_X1 g689(.A(KEYINPUT62), .B(G169gat), .C1(new_n886_), .C2(new_n398_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(G1348gat));
  INV_X1    g691(.A(new_n400_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n886_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n349_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n830_), .A2(new_n885_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(G176gat), .A3(new_n349_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n896_), .A2(new_n899_), .A3(G176gat), .A4(new_n349_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n895_), .B1(new_n898_), .B2(new_n900_), .ZN(G1349gat));
  AOI21_X1  g700(.A(G183gat), .B1(new_n896_), .B2(new_n372_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n886_), .A2(new_n418_), .A3(new_n373_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n886_), .B2(new_n665_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n294_), .A2(new_n567_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n886_), .B2(new_n906_), .ZN(G1351gat));
  NOR2_X1   g706(.A1(new_n696_), .A2(new_n608_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n867_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n398_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n461_), .ZN(G1352gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n628_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n459_), .ZN(G1353gat));
  NAND3_X1  g712(.A1(new_n867_), .A2(new_n372_), .A3(new_n908_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AND2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  OAI21_X1  g717(.A(G218gat), .B1(new_n909_), .B2(new_n665_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n294_), .A2(G218gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n909_), .B2(new_n920_), .ZN(G1355gat));
endmodule


