//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(new_n205_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n207_), .B1(new_n210_), .B2(KEYINPUT85), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n203_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OR3_X1    g020(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(new_n221_), .A3(new_n210_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G71gat), .B(G99gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G43gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n224_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n229_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n227_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G227gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(G15gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n234_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G78gat), .B(G106gat), .ZN(new_n242_));
  INV_X1    g041(.A(G197gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G204gat), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G197gat), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT90), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT21), .B1(new_n244_), .B2(KEYINPUT90), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G211gat), .B(G218gat), .Z(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n244_), .A2(new_n246_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G233gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT89), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(G228gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(G228gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT87), .B1(new_n265_), .B2(KEYINPUT86), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT2), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n266_), .A2(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n269_), .A2(KEYINPUT2), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n269_), .A2(KEYINPUT2), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT86), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(KEYINPUT3), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n277_), .A2(KEYINPUT3), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n267_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(KEYINPUT1), .B2(new_n285_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n285_), .A2(KEYINPUT1), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n273_), .A2(new_n267_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n282_), .A2(new_n286_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n257_), .B(new_n264_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n282_), .A2(new_n286_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n264_), .B1(new_n298_), .B2(new_n257_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n242_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n291_), .A2(new_n292_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G22gat), .B(G50gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT28), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n303_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n298_), .A2(new_n257_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n263_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n242_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n293_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n300_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n311_), .A2(new_n300_), .A3(KEYINPUT91), .A4(new_n306_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT92), .Z(new_n318_));
  AOI22_X1  g117(.A1(new_n249_), .A2(new_n253_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n207_), .B(new_n222_), .C1(new_n210_), .C2(KEYINPUT85), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT94), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n209_), .A2(new_n205_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n206_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT94), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n207_), .A4(new_n222_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n216_), .A2(new_n221_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT93), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT93), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n216_), .A2(new_n221_), .A3(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n321_), .A2(new_n325_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n203_), .B1(new_n322_), .B2(new_n212_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n319_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT20), .B1(new_n224_), .B2(new_n257_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n318_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n224_), .B2(new_n257_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n317_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n330_), .A2(new_n331_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n337_), .C1(new_n338_), .C2(new_n257_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G8gat), .B(G36gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n334_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT96), .B1(new_n231_), .B2(new_n232_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n228_), .A2(new_n229_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT96), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n230_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT97), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n291_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n291_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n233_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT97), .B1(new_n291_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n356_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT98), .B(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n357_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT4), .B(new_n355_), .C1(new_n371_), .C2(new_n359_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n291_), .B2(new_n358_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n362_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n348_), .A2(KEYINPUT95), .B1(new_n370_), .B2(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n334_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n344_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n378_), .A2(new_n379_), .A3(KEYINPUT95), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT99), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(KEYINPUT33), .ZN(new_n382_));
  INV_X1    g181(.A(new_n362_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n361_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n362_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n386_), .B2(new_n369_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n361_), .A2(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n375_), .A2(new_n383_), .ZN(new_n389_));
  AND4_X1   g188(.A1(new_n369_), .A2(new_n388_), .A3(new_n389_), .A4(new_n382_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n377_), .B(new_n380_), .C1(new_n387_), .C2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n369_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n368_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n334_), .A2(new_n339_), .A3(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n332_), .A2(new_n333_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n318_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n336_), .B1(new_n338_), .B2(new_n257_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n397_), .A2(new_n398_), .B1(new_n399_), .B2(new_n317_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n394_), .B(new_n396_), .C1(new_n400_), .C2(new_n395_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n315_), .B1(new_n391_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT27), .B(new_n347_), .C1(new_n400_), .C2(new_n344_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n392_), .A2(new_n393_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(KEYINPUT100), .A4(new_n315_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT100), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n302_), .A2(new_n306_), .B1(new_n311_), .B2(new_n300_), .ZN(new_n410_));
  AND4_X1   g209(.A1(KEYINPUT91), .A2(new_n311_), .A3(new_n300_), .A4(new_n306_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n392_), .B(new_n393_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n404_), .A2(new_n405_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n241_), .B1(new_n402_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT101), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT101), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n418_), .B(new_n241_), .C1(new_n402_), .C2(new_n415_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n315_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n406_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n240_), .A2(new_n407_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(G85gat), .A2(G92gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT67), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n430_), .A3(new_n427_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G99gat), .ZN(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT6), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT8), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n432_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n441_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT68), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n440_), .A2(new_n448_), .A3(new_n441_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n438_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(KEYINPUT69), .A3(new_n432_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT8), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT69), .B1(new_n450_), .B2(new_n432_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n444_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT10), .B(G99gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT64), .B(G92gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT9), .B1(new_n456_), .B2(G85gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(KEYINPUT65), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(KEYINPUT65), .B2(new_n458_), .ZN(new_n461_));
  OAI221_X1 g260(.A(new_n438_), .B1(G106gat), .B2(new_n455_), .C1(new_n457_), .C2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT66), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n455_), .A2(G106gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT66), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n465_), .B(new_n466_), .C1(new_n457_), .C2(new_n461_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT75), .B(KEYINPUT77), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G36gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G29gat), .ZN(new_n472_));
  INV_X1    g271(.A(G29gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G36gat), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n472_), .A2(new_n474_), .A3(KEYINPUT76), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT76), .B1(new_n472_), .B2(new_n474_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G43gat), .B(G50gat), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT76), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n473_), .A2(G36gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n471_), .A2(G29gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n472_), .A2(new_n474_), .A3(KEYINPUT76), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n479_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n470_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n477_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n484_), .A3(new_n479_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n469_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n454_), .A2(new_n468_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n450_), .A2(new_n432_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(KEYINPUT8), .A3(new_n451_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n495_), .A2(new_n444_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n487_), .A2(new_n469_), .A3(new_n488_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n469_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n486_), .A2(KEYINPUT15), .A3(new_n489_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n491_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT34), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT35), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT79), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n505_), .A2(KEYINPUT35), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n491_), .B(new_n511_), .C1(new_n496_), .C2(new_n502_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n508_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G190gat), .B(G218gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT78), .ZN(new_n515_));
  XOR2_X1   g314(.A(G134gat), .B(G162gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(KEYINPUT36), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT36), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(new_n512_), .B2(new_n509_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n513_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n519_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n508_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n425_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n529_), .A2(KEYINPUT104), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT11), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n536_));
  INV_X1    g335(.A(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT70), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n454_), .A2(new_n542_), .A3(new_n468_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n454_), .B2(new_n468_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n532_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT71), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n496_), .B2(new_n542_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n454_), .A2(new_n542_), .A3(new_n468_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n540_), .A2(KEYINPUT72), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n551_), .B(new_n535_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n454_), .B2(new_n468_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n548_), .A2(new_n531_), .A3(new_n549_), .A4(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n557_), .B(new_n532_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n546_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT74), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n546_), .A2(new_n556_), .A3(new_n558_), .A4(new_n563_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G169gat), .B(G197gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT83), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n486_), .A2(KEYINPUT83), .A3(new_n489_), .ZN(new_n579_));
  INV_X1    g378(.A(G1gat), .ZN(new_n580_));
  INV_X1    g379(.A(G8gat), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT14), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G22gat), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n236_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(G15gat), .A2(G22gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT80), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT80), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n582_), .B(new_n588_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G1gat), .B(G8gat), .Z(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n578_), .A2(new_n579_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n578_), .A2(new_n579_), .A3(new_n594_), .A4(KEYINPUT84), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n502_), .A2(new_n594_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n576_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n594_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n603_));
  AOI211_X1 g402(.A(new_n575_), .B(new_n603_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n574_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n603_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n576_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n574_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n600_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n607_), .B(new_n608_), .C1(new_n576_), .C2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n571_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n587_), .A2(new_n589_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n590_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n591_), .ZN(new_n617_));
  AND2_X1   g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n550_), .A2(new_n552_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n620_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n621_), .A2(KEYINPUT17), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT82), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n626_), .B(KEYINPUT17), .Z(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n619_), .B2(new_n542_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n542_), .B2(new_n619_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n529_), .B2(KEYINPUT104), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n530_), .A2(new_n613_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n407_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n425_), .A2(new_n611_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n519_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n524_), .A2(new_n525_), .A3(new_n523_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT37), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n633_), .A3(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n639_), .A2(new_n571_), .A3(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  AOI21_X1  g447(.A(G1gat), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n394_), .A3(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n648_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n638_), .A2(new_n652_), .ZN(G1324gat));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n581_), .A3(new_n413_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n530_), .A2(new_n635_), .A3(new_n613_), .A4(new_n413_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(new_n656_), .A3(G8gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n655_), .B2(G8gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1325gat));
  AOI21_X1  g460(.A(new_n236_), .B1(new_n636_), .B2(new_n240_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n646_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n663_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(G1326gat));
  NAND3_X1  g466(.A1(new_n646_), .A2(new_n583_), .A3(new_n315_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G22gat), .B1(new_n637_), .B2(new_n420_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n613_), .A2(new_n634_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n522_), .A2(new_n526_), .A3(new_n640_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT37), .B1(new_n642_), .B2(new_n643_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT106), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT106), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n675_), .B1(new_n425_), .B2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n678_), .A2(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n423_), .B1(new_n416_), .B2(KEYINPUT101), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n419_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n674_), .B1(new_n682_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n674_), .C1(new_n682_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n407_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n639_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n571_), .A2(new_n528_), .A3(new_n633_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n473_), .A3(new_n394_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n692_), .A2(new_n697_), .ZN(G1328gat));
  NOR2_X1   g497(.A1(new_n406_), .A2(G36gat), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n425_), .A2(new_n611_), .A3(new_n694_), .A4(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT108), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT45), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  INV_X1    g502(.A(new_n690_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n425_), .A2(new_n683_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n685_), .A2(new_n419_), .B1(new_n680_), .B2(new_n679_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n675_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT44), .B1(new_n707_), .B2(new_n674_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n704_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n703_), .B1(new_n709_), .B2(new_n413_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n689_), .A2(new_n703_), .A3(new_n413_), .A4(new_n690_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G36gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n702_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n702_), .B(new_n714_), .C1(new_n710_), .C2(new_n712_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  NAND4_X1  g517(.A1(new_n709_), .A2(KEYINPUT110), .A3(G43gat), .A4(new_n240_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT111), .B(G43gat), .Z(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n695_), .B2(new_n241_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n240_), .A2(G43gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n691_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n721_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT47), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n719_), .A2(new_n724_), .A3(new_n727_), .A4(new_n721_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1330gat));
  AOI21_X1  g528(.A(G50gat), .B1(new_n696_), .B2(new_n315_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n315_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n709_), .B2(new_n731_), .ZN(G1331gat));
  INV_X1    g531(.A(new_n570_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n425_), .A2(new_n612_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(KEYINPUT112), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(KEYINPUT112), .B2(new_n736_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(new_n645_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n407_), .B1(new_n739_), .B2(KEYINPUT113), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(KEYINPUT113), .B2(new_n739_), .ZN(new_n741_));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n735_), .A2(new_n611_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n530_), .A2(new_n635_), .A3(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n407_), .A2(new_n742_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n741_), .A2(new_n742_), .B1(new_n744_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(new_n739_), .ZN(new_n747_));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n413_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n744_), .A2(new_n413_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G64gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT48), .B(new_n748_), .C1(new_n744_), .C2(new_n413_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n747_), .A2(new_n755_), .A3(new_n240_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n744_), .A2(new_n240_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G71gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT49), .B(new_n755_), .C1(new_n744_), .C2(new_n240_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1334gat));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n747_), .A2(new_n762_), .A3(new_n315_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n744_), .A2(new_n315_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(G78gat), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT50), .B(new_n762_), .C1(new_n744_), .C2(new_n315_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1335gat));
  NOR3_X1   g567(.A1(new_n738_), .A2(new_n528_), .A3(new_n633_), .ZN(new_n769_));
  INV_X1    g568(.A(G85gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n394_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n743_), .A2(new_n634_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT114), .Z(new_n773_));
  AND2_X1   g572(.A1(new_n707_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n394_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n770_), .B2(new_n776_), .ZN(G1336gat));
  AOI21_X1  g576(.A(G92gat), .B1(new_n769_), .B2(new_n413_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n413_), .A2(new_n456_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n774_), .B2(new_n779_), .ZN(G1337gat));
  NOR2_X1   g579(.A1(new_n241_), .A2(new_n455_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n769_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n774_), .A2(new_n240_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G99gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g585(.A1(new_n420_), .A2(G106gat), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n773_), .B(new_n315_), .C1(new_n682_), .C2(new_n686_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n788_), .B2(G106gat), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n769_), .A2(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n789_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT52), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  NOR3_X1   g598(.A1(new_n421_), .A2(new_n407_), .A3(new_n241_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n611_), .A2(new_n568_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT117), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n611_), .A2(new_n804_), .A3(new_n568_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n543_), .A2(new_n554_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n531_), .B1(new_n806_), .B2(new_n548_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n556_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n549_), .B1(new_n496_), .B2(new_n553_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n547_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n454_), .A2(new_n468_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n542_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NOR4_X1   g613(.A1(new_n810_), .A2(new_n814_), .A3(new_n808_), .A4(new_n532_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n809_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n565_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n819_), .B(new_n564_), .C1(new_n809_), .C2(new_n816_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n803_), .B(new_n805_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n609_), .A2(new_n576_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n603_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n822_), .B(new_n608_), .C1(new_n823_), .C2(new_n576_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n824_), .A2(new_n605_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n566_), .A2(new_n568_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n527_), .B1(new_n821_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT57), .B1(new_n828_), .B2(KEYINPUT118), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n611_), .A2(new_n804_), .A3(new_n568_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n804_), .B1(new_n611_), .B2(new_n568_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n810_), .A2(new_n814_), .A3(new_n532_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n532_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(KEYINPUT55), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n565_), .B1(new_n837_), .B2(new_n815_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n819_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n565_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n834_), .A2(new_n841_), .B1(new_n826_), .B2(new_n825_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n830_), .B(new_n831_), .C1(new_n842_), .C2(new_n527_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n824_), .A2(new_n605_), .A3(new_n568_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n678_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n841_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n844_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n829_), .A2(new_n843_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n634_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n645_), .A2(new_n571_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n612_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n645_), .A2(new_n571_), .A3(KEYINPUT116), .A4(new_n611_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n678_), .A2(new_n735_), .A3(new_n612_), .A4(new_n633_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT116), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n854_), .A3(new_n612_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n801_), .B1(new_n853_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865_), .B2(new_n611_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT120), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n858_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n861_), .A2(new_n862_), .A3(KEYINPUT54), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n634_), .B2(new_n852_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n869_), .B(KEYINPUT59), .C1(new_n873_), .C2(new_n801_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n868_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n853_), .A2(new_n864_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n867_), .A3(new_n800_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n612_), .A2(KEYINPUT121), .ZN(new_n879_));
  MUX2_X1   g678(.A(KEYINPUT121), .B(new_n879_), .S(G113gat), .Z(new_n880_));
  AOI21_X1  g679(.A(new_n866_), .B1(new_n878_), .B2(new_n880_), .ZN(G1340gat));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n735_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n875_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n735_), .B2(KEYINPUT60), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n882_), .A2(KEYINPUT60), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n876_), .A2(new_n800_), .A3(new_n885_), .A4(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT122), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n884_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n887_), .B(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n877_), .A2(new_n571_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n891_), .B(new_n892_), .C1(new_n894_), .C2(new_n882_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n889_), .A2(new_n895_), .ZN(G1341gat));
  INV_X1    g695(.A(G127gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n865_), .A2(new_n897_), .A3(new_n633_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n875_), .A2(new_n633_), .A3(new_n877_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1342gat));
  AOI21_X1  g699(.A(G134gat), .B1(new_n865_), .B2(new_n527_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT124), .B(G134gat), .Z(new_n902_));
  NOR2_X1   g701(.A1(new_n678_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n878_), .B2(new_n903_), .ZN(G1343gat));
  NOR2_X1   g703(.A1(new_n873_), .A2(new_n240_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n420_), .A2(new_n407_), .A3(new_n413_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n611_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n571_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g711(.A1(new_n907_), .A2(new_n634_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT61), .B(G155gat), .Z(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n908_), .B2(new_n527_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n681_), .A2(G162gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n908_), .B2(new_n917_), .ZN(G1347gat));
  XOR2_X1   g717(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n919_));
  NOR3_X1   g718(.A1(new_n422_), .A2(new_n315_), .A3(new_n406_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n876_), .A2(new_n920_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n921_), .A2(new_n611_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT22), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n919_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G169gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n219_), .B1(new_n922_), .B2(new_n919_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n926_), .ZN(G1348gat));
  NAND2_X1  g726(.A1(new_n921_), .A2(new_n571_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT126), .B(G176gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n921_), .A2(new_n633_), .ZN(new_n931_));
  MUX2_X1   g730(.A(new_n214_), .B(G183gat), .S(new_n931_), .Z(G1350gat));
  NAND3_X1  g731(.A1(new_n921_), .A2(new_n215_), .A3(new_n527_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n678_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n921_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(G190gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n406_), .A2(new_n412_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n905_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n612_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n243_), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n735_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n245_), .ZN(G1353gat));
  INV_X1    g742(.A(new_n939_), .ZN(new_n944_));
  AOI211_X1 g743(.A(KEYINPUT63), .B(G211gat), .C1(new_n944_), .C2(new_n633_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT63), .B(G211gat), .Z(new_n946_));
  AND3_X1   g745(.A1(new_n944_), .A2(new_n633_), .A3(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n944_), .B2(new_n527_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n934_), .A2(G218gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT127), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n944_), .B2(new_n951_), .ZN(G1355gat));
endmodule


