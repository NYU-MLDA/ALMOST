//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  AND2_X1   g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G85gat), .B(G92gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  OAI221_X1 g013(.A(new_n212_), .B1(new_n210_), .B2(new_n213_), .C1(G106gat), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n206_), .A2(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT7), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n213_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n216_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  AOI211_X1 g024(.A(KEYINPUT8), .B(new_n213_), .C1(new_n222_), .C2(new_n219_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n215_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(KEYINPUT11), .B2(new_n228_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT65), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n232_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n204_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n227_), .B(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT12), .A3(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT12), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n240_), .A2(new_n203_), .A3(new_n233_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G120gat), .B(G148gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT5), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G176gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G204gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT67), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n237_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n202_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT68), .B1(new_n244_), .B2(new_n250_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT13), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT13), .B1(new_n253_), .B2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(KEYINPUT69), .A3(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G29gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT71), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G43gat), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n266_), .A2(KEYINPUT71), .ZN(new_n269_));
  INV_X1    g068(.A(G43gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(KEYINPUT71), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n268_), .A2(new_n272_), .A3(G50gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(G50gat), .B1(new_n268_), .B2(new_n272_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n265_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT15), .A3(new_n273_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G22gat), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  INV_X1    g080(.A(G8gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G8gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n279_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G229gat), .A2(G233gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n274_), .A2(new_n275_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n286_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n289_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n291_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n290_), .A2(new_n286_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n264_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n264_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G141gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT78), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n299_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT104), .B1(new_n263_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT104), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n308_), .B(new_n305_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n227_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n239_), .A2(new_n279_), .B1(new_n290_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT72), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G232gat), .A2(G233gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT35), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n316_), .A2(KEYINPUT35), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n313_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n239_), .A2(new_n279_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n311_), .A2(new_n290_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n322_), .A2(KEYINPUT72), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n320_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n322_), .A2(new_n318_), .A3(new_n323_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n324_), .B(new_n325_), .C1(new_n326_), .C2(new_n317_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G190gat), .B(G218gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT73), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G134gat), .ZN(new_n331_));
  INV_X1    g130(.A(G162gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT36), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n333_), .B(KEYINPUT36), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n321_), .A2(new_n327_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT105), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n232_), .B(new_n286_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G231gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G155gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT16), .ZN(new_n346_));
  INV_X1    g145(.A(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G211gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n344_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT76), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n344_), .B(KEYINPUT75), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n351_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n341_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT0), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G57gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(G127gat), .B(G134gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G113gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G120gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  INV_X1    g168(.A(G141gat), .ZN(new_n370_));
  INV_X1    g169(.A(G148gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT83), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT2), .ZN(new_n373_));
  OR3_X1    g172(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT2), .ZN(new_n375_));
  OAI211_X1 g174(.A(KEYINPUT83), .B(new_n375_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT81), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(G155gat), .A3(G162gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n383_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n385_), .B2(KEYINPUT1), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT82), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n381_), .A2(new_n383_), .A3(new_n390_), .A4(new_n387_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G141gat), .B(G148gat), .Z(new_n393_));
  AOI221_X4 g192(.A(new_n369_), .B1(new_n378_), .B2(new_n384_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n378_), .A2(new_n384_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT84), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n368_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT92), .ZN(new_n399_));
  INV_X1    g198(.A(new_n368_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n402_), .B(new_n368_), .C1(new_n394_), .C2(new_n397_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n399_), .A2(KEYINPUT4), .A3(new_n401_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n398_), .A2(KEYINPUT4), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n365_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n399_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n365_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n364_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n399_), .A2(new_n403_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n413_), .A2(new_n405_), .A3(KEYINPUT4), .A4(new_n401_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n404_), .A2(KEYINPUT93), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n407_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n365_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n363_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n412_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G228gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(G233gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(G233gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n303_), .A2(G204gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT86), .B(G204gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n303_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G211gat), .B(G218gat), .Z(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT21), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G197gat), .A2(G204gat), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT21), .B(new_n432_), .C1(new_n427_), .C2(G197gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT87), .ZN(new_n434_));
  INV_X1    g233(.A(G204gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT86), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G204gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n303_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT21), .A4(new_n432_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n429_), .B1(new_n434_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT21), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n426_), .C1(new_n427_), .C2(new_n303_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n431_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n425_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT88), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n425_), .C1(new_n446_), .C2(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n446_), .A2(new_n425_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n394_), .A2(new_n397_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n447_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n458_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n460_), .A3(new_n456_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n397_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n395_), .A2(KEYINPUT84), .A3(new_n396_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n447_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G22gat), .B(G50gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n455_), .A2(new_n447_), .A3(new_n465_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n464_), .A2(new_n466_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n465_), .B1(new_n455_), .B2(new_n447_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n459_), .A2(new_n461_), .A3(new_n471_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n471_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n453_), .A2(new_n460_), .A3(new_n456_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n460_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n483_));
  INV_X1    g282(.A(G169gat), .ZN(new_n484_));
  INV_X1    g283(.A(G176gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(G169gat), .A2(G176gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G183gat), .A2(G190gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT23), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT25), .B(G183gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G190gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n492_), .B(new_n493_), .C1(G183gat), .C2(G190gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G169gat), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n495_), .A2(new_n498_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AOI211_X1 g301(.A(new_n431_), .B(new_n502_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n429_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n444_), .B1(new_n439_), .B2(new_n303_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n441_), .B1(new_n506_), .B2(new_n432_), .ZN(new_n507_));
  AOI21_X1  g306(.A(G197gat), .B1(new_n436_), .B2(new_n438_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n432_), .ZN(new_n509_));
  NOR4_X1   g308(.A1(new_n508_), .A2(KEYINPUT87), .A3(new_n444_), .A4(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n445_), .B(new_n505_), .C1(new_n507_), .C2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n504_), .B1(new_n511_), .B2(new_n430_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT20), .B1(new_n503_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G226gat), .A2(G233gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT90), .Z(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT19), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G64gat), .B(G92gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G8gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(KEYINPUT20), .B(new_n516_), .C1(new_n503_), .C2(new_n512_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n518_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n518_), .B2(new_n524_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n482_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT100), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT100), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n529_), .B(new_n482_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT99), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT99), .B(new_n523_), .C1(new_n518_), .C2(new_n524_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n535_), .B(new_n516_), .C1(new_n503_), .C2(new_n512_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n518_), .A2(new_n524_), .A3(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n513_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n482_), .B1(new_n539_), .B2(new_n523_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n528_), .A2(new_n530_), .B1(new_n534_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n481_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT79), .B(G43gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n502_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(G15gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G71gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n544_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT30), .B(G99gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT80), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n368_), .B(KEYINPUT31), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n420_), .A2(new_n542_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n412_), .A2(new_n419_), .A3(new_n541_), .A4(new_n480_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT101), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n416_), .A2(new_n417_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n363_), .B1(new_n563_), .B2(new_n410_), .ZN(new_n564_));
  AOI211_X1 g363(.A(new_n364_), .B(new_n411_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n528_), .A2(new_n530_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n534_), .A2(new_n540_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n567_), .A2(new_n480_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT101), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n523_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT32), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n518_), .A2(new_n524_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n575_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n574_), .B1(new_n579_), .B2(new_n576_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n412_), .A2(new_n419_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(KEYINPUT33), .B(new_n364_), .C1(new_n408_), .C2(new_n411_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n564_), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n418_), .B2(new_n363_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n525_), .A2(new_n526_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n406_), .A2(KEYINPUT96), .A3(new_n365_), .A4(new_n407_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n363_), .B1(new_n409_), .B2(new_n365_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n589_), .A2(new_n590_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n582_), .B1(new_n587_), .B2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n572_), .B1(new_n599_), .B2(new_n481_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n560_), .B1(new_n600_), .B2(new_n557_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n310_), .A2(new_n359_), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n566_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n305_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n321_), .A2(new_n327_), .A3(new_n338_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n321_), .A2(new_n327_), .B1(new_n334_), .B2(new_n333_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n606_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n358_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n605_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT102), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n605_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n616_), .A2(new_n281_), .A3(new_n420_), .A4(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT103), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(KEYINPUT103), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n603_), .B1(new_n623_), .B2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n541_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n310_), .A2(new_n359_), .A3(new_n626_), .A4(new_n601_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G8gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT39), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n630_), .A3(G8gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n616_), .A2(new_n282_), .A3(new_n626_), .A4(new_n618_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT106), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  INV_X1    g435(.A(new_n631_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n630_), .B1(new_n627_), .B2(G8gat), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n633_), .B(new_n636_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(KEYINPUT40), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  INV_X1    g440(.A(new_n639_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n636_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(G1325gat));
  OAI21_X1  g444(.A(G15gat), .B1(new_n602_), .B2(new_n558_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT41), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n616_), .A2(new_n618_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n557_), .A2(new_n546_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n602_), .B2(new_n481_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n481_), .A2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n648_), .B2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n590_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n412_), .B2(new_n588_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n656_), .A2(new_n585_), .A3(new_n597_), .A4(new_n586_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n480_), .B1(new_n657_), .B2(new_n582_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n558_), .B1(new_n658_), .B2(new_n572_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT43), .B(new_n612_), .C1(new_n659_), .C2(new_n560_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n601_), .B2(new_n613_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n358_), .B(new_n310_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n562_), .A2(new_n571_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT94), .B1(new_n564_), .B2(KEYINPUT33), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n418_), .A2(new_n584_), .A3(new_n588_), .A4(new_n363_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n598_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n581_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n671_), .B2(new_n480_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n559_), .B1(new_n672_), .B2(new_n558_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n673_), .B2(new_n612_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n601_), .A2(new_n661_), .A3(new_n613_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n358_), .A4(new_n310_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n665_), .A2(new_n420_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G29gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n340_), .A2(new_n358_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n601_), .A2(new_n604_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n566_), .A2(G29gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n682_), .A2(new_n686_), .A3(new_n626_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n688_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n682_), .A2(new_n686_), .A3(new_n626_), .A4(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n665_), .A2(new_n626_), .A3(new_n677_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G36gat), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n694_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n665_), .A2(new_n557_), .A3(new_n677_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G43gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n682_), .A2(new_n270_), .A3(new_n557_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1330gat));
  AND3_X1   g506(.A1(new_n665_), .A2(new_n480_), .A3(new_n677_), .ZN(new_n708_));
  INV_X1    g507(.A(G50gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n480_), .A2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT110), .Z(new_n711_));
  OAI22_X1  g510(.A1(new_n708_), .A2(new_n709_), .B1(new_n683_), .B2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n263_), .A2(new_n306_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n601_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n359_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n566_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n614_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n420_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n716_), .B2(new_n720_), .ZN(G1332gat));
  OAI21_X1  g520(.A(G64gat), .B1(new_n715_), .B2(new_n541_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT48), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n541_), .A2(G64gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT111), .Z(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n718_), .B2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n715_), .B2(new_n558_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n548_), .A3(new_n557_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n715_), .B2(new_n481_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n481_), .A2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n718_), .B2(new_n733_), .ZN(G1335gat));
  NAND2_X1  g533(.A1(new_n714_), .A2(new_n681_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n420_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n676_), .A2(new_n358_), .A3(new_n713_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n420_), .A2(G85gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n736_), .B2(new_n626_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n626_), .A2(G92gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n739_), .B2(new_n743_), .ZN(G1337gat));
  NAND4_X1  g543(.A1(new_n676_), .A2(new_n358_), .A3(new_n557_), .A4(new_n713_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n745_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT112), .B1(new_n745_), .B2(G99gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n735_), .A2(new_n214_), .A3(new_n558_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(KEYINPUT51), .A4(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(G99gat), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n745_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n750_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n751_), .A2(new_n759_), .ZN(G1338gat));
  OR3_X1    g559(.A1(new_n735_), .A2(G106gat), .A3(new_n481_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n676_), .A2(new_n358_), .A3(new_n480_), .A4(new_n713_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g566(.A1(new_n566_), .A2(new_n542_), .A3(new_n558_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n243_), .A2(KEYINPUT117), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n240_), .A2(new_n242_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n204_), .B1(new_n772_), .B2(new_n234_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT117), .B1(new_n243_), .B2(new_n770_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  XOR2_X1   g574(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n243_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n243_), .A2(new_n779_), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n250_), .B1(new_n775_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n250_), .C1(new_n775_), .C2(new_n781_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n783_), .A2(new_n306_), .A3(new_n252_), .A4(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n297_), .A2(new_n298_), .A3(new_n304_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n288_), .A2(new_n293_), .A3(new_n291_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n289_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n304_), .ZN(new_n791_));
  OR3_X1    g590(.A1(new_n787_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n787_), .B2(new_n791_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n254_), .B2(new_n253_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n340_), .B1(new_n786_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n783_), .A2(new_n252_), .A3(new_n794_), .A4(new_n785_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n802_), .B2(new_n613_), .ZN(new_n803_));
  AOI211_X1 g602(.A(KEYINPUT119), .B(new_n612_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n800_), .A2(new_n801_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n798_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n802_), .A2(new_n613_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT119), .ZN(new_n810_));
  INV_X1    g609(.A(new_n805_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n802_), .A2(new_n799_), .A3(new_n613_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT120), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n358_), .B1(new_n808_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n358_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n612_), .A2(new_n816_), .A3(new_n305_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n259_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT114), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n817_), .A2(new_n818_), .A3(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(KEYINPUT54), .C1(new_n817_), .C2(new_n818_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n769_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825_), .B2(new_n306_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n786_), .A2(new_n795_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n340_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n797_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n813_), .B2(KEYINPUT120), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n806_), .A2(new_n807_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n816_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n824_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT59), .B(new_n768_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n769_), .A2(KEYINPUT121), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n769_), .A2(KEYINPUT121), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n816_), .B1(new_n813_), .B2(new_n798_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n839_), .C1(new_n840_), .C2(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n305_), .B1(new_n837_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n826_), .B1(new_n844_), .B2(G113gat), .ZN(G1340gat));
  AOI21_X1  g644(.A(new_n263_), .B1(new_n837_), .B2(new_n843_), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n825_), .B1(KEYINPUT60), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n263_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n850_));
  AOI21_X1  g649(.A(G120gat), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n846_), .A2(new_n847_), .B1(new_n848_), .B2(new_n851_), .ZN(G1341gat));
  NAND2_X1  g651(.A1(new_n816_), .A2(G127gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT122), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n837_), .B2(new_n843_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n825_), .A2(new_n816_), .ZN(new_n858_));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G127gat), .B1(new_n825_), .B2(new_n816_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT123), .B1(new_n856_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n825_), .B2(new_n341_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n612_), .B1(new_n837_), .B2(new_n843_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT124), .B(G134gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n481_), .A2(new_n557_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n566_), .A2(new_n626_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n370_), .A3(new_n306_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G141gat), .B1(new_n874_), .B2(new_n305_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n371_), .A3(new_n849_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G148gat), .B1(new_n874_), .B2(new_n263_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1345gat));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n875_), .B2(new_n816_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n883_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n874_), .A2(new_n358_), .A3(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1346gat));
  NOR3_X1   g686(.A1(new_n874_), .A2(new_n332_), .A3(new_n612_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n875_), .A2(new_n341_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n332_), .B2(new_n889_), .ZN(G1347gat));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n420_), .A2(new_n558_), .A3(new_n541_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n481_), .B(new_n892_), .C1(new_n840_), .C2(new_n836_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n305_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT22), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n484_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n891_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G169gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n896_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(G1348gat));
  INV_X1    g700(.A(new_n893_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902_), .B2(new_n849_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n480_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n849_), .A2(G176gat), .A3(new_n892_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NOR3_X1   g705(.A1(new_n893_), .A2(new_n358_), .A3(new_n496_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n816_), .A3(new_n892_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n347_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n902_), .A2(new_n341_), .A3(new_n497_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G190gat), .B1(new_n893_), .B2(new_n612_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  NOR2_X1   g711(.A1(new_n871_), .A2(new_n420_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n541_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n917_), .B(new_n918_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n305_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n303_), .ZN(G1352gat));
  OAI21_X1  g720(.A(G204gat), .B1(new_n919_), .B2(new_n263_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n916_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n923_), .A2(new_n849_), .A3(new_n439_), .A4(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT127), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n922_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1353gat));
  INV_X1    g728(.A(new_n919_), .ZN(new_n930_));
  AOI211_X1 g729(.A(KEYINPUT63), .B(G211gat), .C1(new_n930_), .C2(new_n816_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT63), .B(G211gat), .Z(new_n932_));
  AND3_X1   g731(.A1(new_n930_), .A2(new_n816_), .A3(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1354gat));
  INV_X1    g733(.A(G218gat), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n919_), .A2(new_n935_), .A3(new_n612_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n930_), .A2(new_n341_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n935_), .ZN(G1355gat));
endmodule


