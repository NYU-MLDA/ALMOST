//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G183gat), .B(G211gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT86), .B1(new_n206_), .B2(KEYINPUT17), .ZN(new_n207_));
  AND2_X1   g006(.A1(G231gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G1gat), .A2(G8gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT14), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G15gat), .A2(G22gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(G15gat), .A2(G22gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT84), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT84), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n211_), .B(new_n216_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G1gat), .B(G8gat), .Z(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n215_), .A2(new_n219_), .A3(new_n217_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n209_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n209_), .A2(new_n224_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G78gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT70), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n230_), .B2(KEYINPUT11), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(KEYINPUT70), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n229_), .A2(KEYINPUT70), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(KEYINPUT11), .A3(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239_));
  INV_X1    g038(.A(new_n206_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n227_), .A2(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n225_), .A2(new_n237_), .A3(new_n226_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G190gat), .B(G218gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(G134gat), .B(G162gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT36), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT82), .Z(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT65), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT6), .ZN(new_n256_));
  AND2_X1   g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n252_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n257_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n255_), .A2(KEYINPUT6), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n253_), .A2(KEYINPUT65), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(KEYINPUT66), .A3(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT64), .B(G85gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT9), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(G92gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n272_));
  INV_X1    g071(.A(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(G85gat), .A2(G92gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G85gat), .A2(G92gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT9), .A3(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n260_), .A2(new_n266_), .A3(new_n271_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT71), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n278_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(new_n270_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n260_), .A4(new_n266_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(G85gat), .A2(G92gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G85gat), .A2(G92gat), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n287_), .A2(new_n288_), .A3(KEYINPUT68), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n264_), .A2(new_n265_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT7), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G99gat), .A2(G106gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n292_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n292_), .B(KEYINPUT69), .C1(new_n293_), .C2(new_n299_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT8), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n299_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n260_), .A2(new_n305_), .A3(new_n266_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n289_), .A2(new_n291_), .A3(KEYINPUT8), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n286_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT15), .ZN(new_n310_));
  XOR2_X1   g109(.A(G29gat), .B(G36gat), .Z(new_n311_));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G29gat), .B(G36gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT77), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G43gat), .B(G50gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n310_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n315_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n316_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT15), .A3(new_n317_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT78), .B1(new_n309_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n286_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n303_), .A2(KEYINPUT8), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT7), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT67), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n296_), .B1(new_n295_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n332_), .A2(new_n264_), .A3(new_n265_), .A4(new_n297_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT69), .B1(new_n333_), .B2(new_n292_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n308_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337_));
  INV_X1    g136(.A(new_n325_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n326_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G232gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT76), .B(KEYINPUT35), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n343_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n344_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n323_), .A2(new_n317_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n335_), .A2(new_n280_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT79), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n335_), .A2(new_n353_), .A3(new_n280_), .A4(new_n350_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n349_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n340_), .A2(new_n346_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n346_), .B1(new_n340_), .B2(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n251_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n337_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n359_));
  AOI211_X1 g158(.A(KEYINPUT78), .B(new_n325_), .C1(new_n327_), .C2(new_n335_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n349_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n280_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n353_), .B1(new_n364_), .B2(new_n350_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n354_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n345_), .B1(new_n361_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n340_), .A2(new_n355_), .A3(new_n346_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT36), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n249_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n358_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(KEYINPUT37), .ZN(new_n377_));
  INV_X1    g176(.A(new_n250_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT37), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n358_), .B2(new_n374_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n376_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n246_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  NOR3_X1   g187(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT23), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G183gat), .A3(G190gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n389_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G190gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n394_), .B(new_n397_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G183gat), .ZN(new_n403_));
  INV_X1    g202(.A(G190gat), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n391_), .A2(new_n393_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT94), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G169gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n405_), .B2(KEYINPUT94), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n402_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT99), .ZN(new_n411_));
  AND2_X1   g210(.A1(G197gat), .A2(G204gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G197gat), .A2(G204gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G211gat), .B(G218gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n412_), .A2(new_n413_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT21), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT100), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT21), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G211gat), .B(G218gat), .Z(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n413_), .B2(new_n412_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n421_), .B1(new_n425_), .B2(new_n416_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n422_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT100), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n410_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n419_), .A2(new_n422_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n405_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n408_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n402_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT20), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n388_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G8gat), .B(G36gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT18), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n423_), .A2(new_n428_), .A3(new_n410_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n388_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n435_), .A2(new_n439_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT105), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n429_), .A2(new_n434_), .A3(new_n388_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n442_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n388_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n439_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n447_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT105), .B(new_n439_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT27), .B(new_n446_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n439_), .B1(new_n435_), .B2(new_n444_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n445_), .A2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(KEYINPUT27), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(G85gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT0), .B(G57gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  XOR2_X1   g265(.A(G127gat), .B(G134gat), .Z(new_n467_));
  XOR2_X1   g266(.A(G113gat), .B(G120gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT96), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G134gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G120gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT95), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G155gat), .A2(G162gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G141gat), .A2(G148gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT3), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n486_), .B1(G141gat), .B2(G148gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT97), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT97), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n481_), .B1(KEYINPUT1), .B2(new_n479_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(KEYINPUT1), .B2(new_n479_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G141gat), .B(G148gat), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n473_), .B(new_n478_), .C1(new_n496_), .C2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n488_), .A2(KEYINPUT97), .A3(new_n491_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT97), .B1(new_n488_), .B2(new_n491_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n482_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n469_), .A2(new_n476_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n500_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n466_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n473_), .A2(new_n478_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n500_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT4), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n465_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n502_), .A2(new_n464_), .A3(new_n507_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT102), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT102), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n502_), .A2(new_n516_), .A3(new_n464_), .A4(new_n507_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n463_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n463_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n512_), .A2(new_n520_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n510_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT28), .B1(new_n510_), .B2(KEYINPUT29), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n526_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n430_), .B1(new_n510_), .B2(KEYINPUT29), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G228gat), .A2(G233gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT98), .Z(new_n533_));
  OR2_X1    g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT101), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n510_), .A2(KEYINPUT29), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n538_), .A2(new_n423_), .A3(new_n428_), .A4(new_n533_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n530_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n536_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(new_n529_), .A3(new_n527_), .A4(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G227gat), .A2(G233gat), .ZN(new_n548_));
  INV_X1    g347(.A(G15gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT30), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n410_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(new_n509_), .Z(new_n553_));
  XNOR2_X1  g352(.A(G71gat), .B(G99gat), .ZN(new_n554_));
  INV_X1    g353(.A(G43gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT31), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n553_), .B(new_n557_), .ZN(new_n558_));
  NOR4_X1   g357(.A1(new_n459_), .A2(new_n522_), .A3(new_n547_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n522_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n455_), .A2(new_n560_), .A3(new_n547_), .A4(new_n458_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n439_), .A2(KEYINPUT32), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n429_), .A2(new_n434_), .A3(new_n388_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n443_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n562_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n435_), .A3(new_n444_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n515_), .A2(new_n517_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(KEYINPUT33), .A3(new_n520_), .A4(new_n512_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n464_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n502_), .A2(new_n465_), .A3(new_n507_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n463_), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n457_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT104), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT103), .B(KEYINPUT33), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n521_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n521_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n569_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n561_), .B1(new_n581_), .B2(new_n547_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n559_), .B1(new_n582_), .B2(new_n558_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n364_), .B2(new_n237_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT12), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n336_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n335_), .A2(new_n237_), .A3(new_n280_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n589_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n364_), .A2(new_n237_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n590_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G120gat), .B(G148gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT73), .ZN(new_n597_));
  XOR2_X1   g396(.A(G176gat), .B(G204gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n591_), .A2(new_n595_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n591_), .A2(new_n595_), .A3(new_n604_), .A4(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n591_), .A2(new_n595_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n601_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(KEYINPUT13), .A3(new_n609_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n318_), .A2(new_n319_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n223_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n350_), .A2(new_n222_), .A3(new_n221_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(KEYINPUT88), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT88), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n223_), .A3(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n617_), .A2(G229gat), .A3(G233gat), .A4(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n320_), .A2(new_n223_), .A3(new_n324_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT89), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n616_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT90), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n620_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT91), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n625_), .B1(new_n620_), .B2(new_n624_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT92), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n626_), .A4(new_n630_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n620_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT93), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT93), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n620_), .A2(new_n624_), .A3(new_n639_), .A4(new_n629_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n633_), .A2(new_n636_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n612_), .A2(new_n613_), .A3(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n386_), .A2(new_n583_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n645_), .A2(G1gat), .A3(new_n560_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n246_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n373_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n356_), .A2(new_n357_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n379_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n583_), .A2(new_n649_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n643_), .A2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n612_), .A2(KEYINPUT106), .A3(new_n613_), .A4(new_n642_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n560_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n646_), .A2(new_n647_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n648_), .A2(new_n659_), .A3(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(G8gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n644_), .A2(new_n662_), .A3(new_n459_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  INV_X1    g463(.A(new_n658_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n459_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(G8gat), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT39), .B(new_n662_), .C1(new_n665_), .C2(new_n459_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT40), .B(new_n663_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(new_n558_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n644_), .A2(new_n549_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G15gat), .B1(new_n658_), .B2(new_n558_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n676_), .A2(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(new_n547_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n645_), .A2(G22gat), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G22gat), .B1(new_n658_), .B2(new_n681_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n376_), .A2(new_n384_), .B1(new_n652_), .B2(new_n381_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n375_), .A2(KEYINPUT37), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT83), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n583_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n521_), .A2(new_n577_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT104), .ZN(new_n694_));
  INV_X1    g493(.A(new_n456_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n446_), .A2(new_n574_), .A3(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n694_), .A2(new_n696_), .A3(new_n580_), .A4(new_n571_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n569_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n547_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n560_), .A2(new_n455_), .A3(new_n547_), .A4(new_n458_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n558_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n459_), .A2(new_n547_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n560_), .A3(new_n674_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n383_), .A2(new_n385_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT43), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n692_), .A2(new_n649_), .A3(new_n706_), .A4(new_n657_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n704_), .A2(new_n705_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n246_), .B1(new_n710_), .B2(new_n687_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n711_), .A2(KEYINPUT44), .A3(new_n657_), .A4(new_n706_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(G29gat), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n560_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n652_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n246_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT107), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n583_), .A2(new_n643_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n522_), .A3(new_n719_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n713_), .A2(new_n715_), .B1(new_n714_), .B2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(new_n459_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n719_), .A3(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT45), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n709_), .A2(new_n712_), .A3(new_n459_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G36gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n725_), .B(new_n727_), .C1(KEYINPUT108), .C2(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1329gat));
  NOR2_X1   g531(.A1(new_n558_), .A2(new_n555_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n709_), .A2(new_n712_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT109), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n709_), .A2(new_n712_), .A3(new_n736_), .A4(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n718_), .A2(new_n719_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n555_), .B1(new_n738_), .B2(new_n558_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT47), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n735_), .A2(new_n742_), .A3(new_n737_), .A4(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  NAND4_X1  g543(.A1(new_n709_), .A2(new_n712_), .A3(G50gat), .A4(new_n547_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n738_), .A2(new_n681_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(G50gat), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n612_), .A2(new_n613_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n583_), .A2(new_n751_), .A3(new_n642_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n649_), .A2(new_n652_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n522_), .A2(G57gat), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n386_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n752_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n560_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n757_), .B(new_n758_), .C1(G57gat), .C2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT112), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n754_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n459_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n766_), .A2(new_n767_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n459_), .A2(new_n764_), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n768_), .A2(new_n769_), .B1(new_n760_), .B2(new_n770_), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n754_), .B2(new_n558_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT49), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n558_), .A2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n760_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n754_), .B2(new_n681_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT50), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n681_), .A2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n760_), .B2(new_n778_), .ZN(G1335gat));
  NAND2_X1  g578(.A1(new_n718_), .A2(new_n752_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n522_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n751_), .A2(new_n642_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n711_), .A2(new_n706_), .A3(new_n783_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n784_), .A2(new_n267_), .A3(new_n560_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n782_), .A2(new_n785_), .ZN(G1336gat));
  OAI21_X1  g585(.A(G92gat), .B1(new_n784_), .B2(new_n722_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n722_), .A2(G92gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n780_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n784_), .B2(new_n558_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n674_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n780_), .B2(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n781_), .A2(new_n273_), .A3(new_n547_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n711_), .A2(new_n547_), .A3(new_n706_), .A4(new_n783_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n797_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n797_), .B(new_n805_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n617_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n623_), .B1(new_n224_), .B2(new_n350_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n629_), .B1(new_n810_), .B2(new_n621_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n641_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n590_), .B1(new_n309_), .B2(new_n586_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n335_), .A2(new_n280_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT12), .B1(new_n816_), .B2(new_n238_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n592_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT55), .A3(new_n591_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n815_), .A2(new_n817_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n589_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n608_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n601_), .A2(new_n824_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n819_), .A2(new_n822_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT116), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n819_), .A2(new_n822_), .A3(new_n829_), .A4(new_n826_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n642_), .A2(new_n606_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n814_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n808_), .B1(new_n833_), .B2(new_n652_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n642_), .A2(new_n606_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(KEYINPUT116), .A2(new_n827_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n830_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT57), .B(new_n716_), .C1(new_n837_), .C2(new_n814_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n819_), .A2(new_n822_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n840_), .A2(new_n826_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n606_), .A2(new_n641_), .A3(new_n812_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n825_), .A2(new_n827_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n813_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(KEYINPUT58), .A3(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n688_), .A2(new_n843_), .A3(new_n690_), .A4(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n834_), .A2(new_n838_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n649_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n642_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n612_), .A2(new_n613_), .A3(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT54), .B1(new_n386_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n691_), .A2(new_n853_), .A3(new_n854_), .A4(new_n246_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n849_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n702_), .A2(new_n522_), .A3(new_n674_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(KEYINPUT118), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n834_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT117), .B(new_n808_), .C1(new_n833_), .C2(new_n652_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n838_), .A4(new_n847_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n867_), .A2(new_n649_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n858_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n642_), .B(new_n863_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G113gat), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n867_), .A2(new_n649_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n856_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n859_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  OR3_X1    g674(.A1(new_n875_), .A2(G113gat), .A3(new_n850_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n876_), .ZN(G1340gat));
  OAI211_X1 g676(.A(new_n750_), .B(new_n863_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G120gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT119), .B1(new_n880_), .B2(G120gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(G120gat), .B1(new_n750_), .B2(new_n880_), .ZN(new_n882_));
  MUX2_X1   g681(.A(new_n881_), .B(KEYINPUT119), .S(new_n882_), .Z(new_n883_));
  NAND2_X1  g682(.A1(new_n869_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n884_), .ZN(G1341gat));
  AOI21_X1  g684(.A(G127gat), .B1(new_n869_), .B2(new_n246_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n863_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n875_), .B2(KEYINPUT59), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n649_), .A2(KEYINPUT120), .ZN(new_n889_));
  MUX2_X1   g688(.A(KEYINPUT120), .B(new_n889_), .S(G127gat), .Z(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n888_), .B2(new_n890_), .ZN(G1342gat));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892_));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n892_), .B(new_n893_), .C1(new_n875_), .C2(new_n716_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n868_), .A2(new_n716_), .A3(new_n858_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT121), .B1(new_n895_), .B2(G134gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT122), .B(G134gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n691_), .A2(new_n897_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n894_), .A2(new_n896_), .B1(new_n888_), .B2(new_n898_), .ZN(G1343gat));
  INV_X1    g698(.A(new_n868_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n681_), .A2(new_n674_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n722_), .A2(new_n901_), .A3(new_n522_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(new_n642_), .A3(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g704(.A1(new_n900_), .A2(new_n750_), .A3(new_n903_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g706(.A1(new_n900_), .A2(new_n246_), .A3(new_n903_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  INV_X1    g709(.A(G162gat), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n868_), .A2(new_n911_), .A3(new_n691_), .A4(new_n902_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n900_), .A2(new_n652_), .A3(new_n903_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(KEYINPUT123), .A3(new_n911_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n868_), .A2(new_n716_), .A3(new_n902_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(G162gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n912_), .B1(new_n914_), .B2(new_n917_), .ZN(G1347gat));
  INV_X1    g717(.A(KEYINPUT22), .ZN(new_n919_));
  NOR4_X1   g718(.A1(new_n722_), .A2(new_n522_), .A3(new_n547_), .A4(new_n558_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n642_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n857_), .A2(new_n919_), .A3(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(KEYINPUT62), .A3(new_n398_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n857_), .A2(new_n925_), .A3(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G169gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n921_), .B1(new_n849_), .B2(new_n856_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n928_), .B2(new_n919_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n924_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT124), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n924_), .B(new_n932_), .C1(new_n927_), .C2(new_n929_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1348gat));
  NAND2_X1  g733(.A1(new_n857_), .A2(new_n920_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(G176gat), .B1(new_n936_), .B2(new_n750_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n900_), .A2(new_n920_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n751_), .A2(new_n399_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(G1349gat));
  NOR3_X1   g739(.A1(new_n935_), .A2(new_n649_), .A3(new_n395_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n246_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n403_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n935_), .B2(new_n691_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n396_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n935_), .A2(new_n716_), .A3(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(KEYINPUT125), .B1(new_n945_), .B2(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n947_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n949_), .A2(new_n950_), .A3(new_n944_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n948_), .A2(new_n951_), .ZN(G1351gat));
  NAND3_X1  g751(.A1(new_n901_), .A2(new_n560_), .A3(new_n459_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n868_), .A2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n642_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n750_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g757(.A(new_n649_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n954_), .A2(new_n959_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n960_), .B(new_n963_), .ZN(G1354gat));
  INV_X1    g763(.A(new_n954_), .ZN(new_n965_));
  OAI21_X1  g764(.A(G218gat), .B1(new_n965_), .B2(new_n691_), .ZN(new_n966_));
  INV_X1    g765(.A(G218gat), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n954_), .A2(new_n967_), .A3(new_n652_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1355gat));
endmodule


