//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G127gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G134gat), .ZN(new_n208_));
  INV_X1    g007(.A(G134gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G127gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT83), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n203_), .B1(new_n206_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n204_), .A2(new_n205_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT83), .B1(new_n208_), .B2(new_n210_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n202_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT31), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT84), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT22), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT22), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G169gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT78), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT78), .B1(new_n225_), .B2(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(G176gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT79), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(G176gat), .B1(new_n224_), .B2(KEYINPUT78), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G169gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n232_), .B(new_n233_), .C1(KEYINPUT78), .C2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n239_), .A2(new_n240_), .B1(G169gat), .B2(G176gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n231_), .A2(new_n235_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT25), .B(G183gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT26), .B(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n237_), .A2(G183gat), .A3(G190gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n247_), .A2(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n246_), .B(new_n251_), .C1(new_n250_), .C2(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n242_), .A2(new_n243_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n243_), .B1(new_n242_), .B2(new_n254_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT30), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n242_), .A2(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT80), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(new_n243_), .A3(new_n254_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n258_), .A2(new_n264_), .A3(KEYINPUT81), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(G43gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(G15gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n271_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n268_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n222_), .B1(new_n279_), .B2(new_n218_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n221_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT85), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n284_));
  INV_X1    g083(.A(new_n218_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n283_), .B(new_n284_), .C1(new_n286_), .C2(new_n222_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G228gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT89), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G22gat), .B(G50gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT1), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G155gat), .A3(G162gat), .ZN(new_n300_));
  OR2_X1    g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G141gat), .B(G148gat), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  OR3_X1    g106(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  INV_X1    g108(.A(G141gat), .ZN(new_n310_));
  INV_X1    g109(.A(G148gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n308_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n301_), .A2(new_n297_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n305_), .A2(new_n307_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n296_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G197gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT90), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G197gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n323_), .A3(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT91), .ZN(new_n325_));
  INV_X1    g124(.A(G204gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(G197gat), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT21), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT92), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT92), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n324_), .A2(new_n329_), .A3(new_n333_), .A4(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT91), .B(G204gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT90), .B(G197gat), .ZN(new_n339_));
  OAI22_X1  g138(.A1(new_n338_), .A2(G197gat), .B1(new_n339_), .B2(G204gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n340_), .B2(KEYINPUT21), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT93), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n324_), .A2(new_n329_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n336_), .A2(new_n330_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n324_), .A2(new_n329_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n335_), .A2(new_n341_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(G78gat), .B1(new_n319_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n335_), .A2(new_n341_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n347_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n315_), .A2(new_n316_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n306_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n356_), .A2(KEYINPUT29), .B1(new_n291_), .B2(new_n290_), .ZN(new_n357_));
  INV_X1    g156(.A(G78gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n352_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n349_), .A2(G106gat), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(G106gat), .B1(new_n349_), .B2(new_n359_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n317_), .A2(new_n363_), .A3(new_n318_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT87), .B1(new_n356_), .B2(KEYINPUT29), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n361_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G106gat), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n319_), .A2(new_n348_), .A3(G78gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n358_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n374_), .B1(new_n378_), .B2(new_n360_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n295_), .B1(new_n371_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n370_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n374_), .A3(new_n360_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n294_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n305_), .A2(new_n307_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(new_n353_), .A3(new_n215_), .A4(new_n212_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n216_), .A2(new_n356_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT4), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT101), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(KEYINPUT102), .Z(new_n392_));
  NAND4_X1  g191(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT101), .A4(KEYINPUT4), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n387_), .A2(KEYINPUT4), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT33), .A4(new_n401_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n390_), .A2(new_n391_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n386_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT103), .A3(new_n400_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n400_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT103), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n408_), .A3(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n404_), .A2(new_n405_), .A3(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G8gat), .B(G36gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT19), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n251_), .B(KEYINPUT96), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n253_), .A2(KEYINPUT95), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n250_), .B1(new_n253_), .B2(KEYINPUT95), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n424_), .A2(new_n425_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n239_), .A2(new_n240_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n234_), .A2(new_n229_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n252_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT97), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT97), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n427_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT20), .B(new_n422_), .C1(new_n435_), .C2(new_n352_), .ZN(new_n436_));
  AOI21_X1  g235(.A(G204gat), .B1(new_n321_), .B2(new_n323_), .ZN(new_n437_));
  AOI21_X1  g236(.A(G197gat), .B1(new_n327_), .B2(new_n328_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT21), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n336_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n347_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n255_), .A2(new_n256_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT98), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n262_), .A2(new_n445_), .A3(new_n352_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n257_), .A2(new_n348_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(new_n435_), .B2(new_n352_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n422_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n419_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n435_), .A2(new_n352_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n422_), .A2(KEYINPUT20), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n443_), .A2(KEYINPUT98), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n445_), .B1(new_n262_), .B2(new_n352_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(new_n450_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n421_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n460_), .A3(new_n418_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT100), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n452_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n452_), .B2(new_n461_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n413_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n395_), .A2(new_n396_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n400_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n447_), .A2(new_n451_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n467_), .A2(new_n402_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n448_), .A2(new_n450_), .A3(new_n422_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n348_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT20), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n471_), .B1(new_n474_), .B2(new_n422_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT104), .ZN(new_n476_));
  INV_X1    g275(.A(new_n469_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n470_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n384_), .B1(new_n465_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n471_), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT20), .B(new_n472_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n421_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n418_), .B(KEYINPUT105), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT27), .B(new_n461_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n452_), .A2(new_n461_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT27), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n467_), .A2(new_n402_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n288_), .B1(new_n481_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n380_), .A2(new_n383_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT106), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n283_), .B1(new_n286_), .B2(new_n222_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n486_), .A3(new_n489_), .A4(KEYINPUT106), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n498_), .A2(new_n491_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT71), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n505_), .A2(KEYINPUT71), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n504_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n505_), .A2(KEYINPUT71), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(new_n506_), .A3(new_n503_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515_));
  INV_X1    g314(.A(G1gat), .ZN(new_n516_));
  INV_X1    g315(.A(G8gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G1gat), .B(G8gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n509_), .A2(KEYINPUT15), .A3(new_n511_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n514_), .A2(KEYINPUT77), .A3(new_n522_), .A4(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT76), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n512_), .B2(new_n521_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n512_), .A2(new_n521_), .A3(new_n531_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n530_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n534_), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n537_), .A2(new_n532_), .B1(new_n521_), .B2(new_n512_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n530_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n502_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT65), .ZN(new_n549_));
  INV_X1    g348(.A(G99gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n375_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT7), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(G99gat), .A3(G106gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT7), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n549_), .A2(new_n558_), .A3(new_n550_), .A4(new_n375_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(KEYINPUT8), .A3(new_n563_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT10), .B(G99gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT64), .B(G106gat), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n568_), .A2(new_n569_), .B1(new_n563_), .B2(KEYINPUT9), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n561_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n557_), .A3(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n567_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n566_), .A2(KEYINPUT66), .A3(new_n573_), .A4(new_n567_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(new_n523_), .A3(new_n514_), .A4(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n566_), .A2(new_n567_), .A3(new_n573_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n512_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT70), .Z(new_n585_));
  AND3_X1   g384(.A1(new_n578_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT36), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n586_), .A2(new_n587_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n590_), .B(KEYINPUT36), .Z(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NOR4_X1   g399(.A1(new_n586_), .A2(new_n587_), .A3(new_n600_), .A4(new_n592_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n593_), .A2(KEYINPUT72), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n595_), .B(KEYINPUT73), .Z(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n601_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n599_), .B1(new_n605_), .B2(new_n598_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT11), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT11), .ZN(new_n609_));
  XOR2_X1   g408(.A(G71gat), .B(G78gat), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n521_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n616_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n616_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT74), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n606_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT75), .ZN(new_n629_));
  INV_X1    g428(.A(new_n613_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT12), .B1(new_n574_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n574_), .A2(new_n630_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n611_), .A2(KEYINPUT12), .A3(new_n612_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n576_), .A2(new_n577_), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n634_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n632_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n574_), .A2(new_n630_), .ZN(new_n640_));
  OAI211_X1 g439(.A(G230gat), .B(G233gat), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT5), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n641_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT68), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT68), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n638_), .A2(new_n641_), .A3(new_n648_), .A4(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT67), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n638_), .A2(new_n641_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n645_), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n650_), .A2(new_n654_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n655_));
  INV_X1    g454(.A(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n638_), .A2(new_n641_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n645_), .B1(new_n657_), .B2(KEYINPUT67), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n656_), .A2(new_n658_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n548_), .A2(new_n629_), .A3(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n491_), .A2(G1gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(KEYINPUT38), .A3(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n597_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n494_), .B2(new_n501_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n547_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n663_), .A2(new_n672_), .A3(new_n626_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n491_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n668_), .A2(new_n669_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT107), .ZN(G1324gat));
  NAND3_X1  g476(.A1(new_n664_), .A2(new_n517_), .A3(new_n490_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n490_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G8gat), .B1(new_n674_), .B2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n674_), .B2(new_n288_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT109), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n288_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n664_), .A2(new_n273_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n687_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n690_), .A3(new_n691_), .ZN(G1326gat));
  OAI21_X1  g491(.A(G22gat), .B1(new_n674_), .B2(new_n495_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT42), .ZN(new_n694_));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n664_), .A2(new_n695_), .A3(new_n384_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n627_), .A2(new_n670_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n548_), .A2(new_n663_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n491_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n662_), .A2(new_n547_), .A3(new_n627_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT110), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n606_), .B2(KEYINPUT111), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n502_), .B2(new_n606_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n606_), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n708_), .B(new_n705_), .C1(new_n494_), .C2(new_n501_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n703_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n703_), .B(KEYINPUT44), .C1(new_n707_), .C2(new_n709_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n700_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n701_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n490_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n699_), .A2(new_n719_), .A3(new_n490_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT45), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n699_), .A2(new_n722_), .A3(new_n719_), .A4(new_n490_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n718_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NAND4_X1  g529(.A1(new_n712_), .A2(G43gat), .A3(new_n499_), .A4(new_n713_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n699_), .A2(new_n689_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n270_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n699_), .B2(new_n384_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n384_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n714_), .B2(new_n737_), .ZN(G1331gat));
  NOR3_X1   g537(.A1(new_n662_), .A2(new_n547_), .A3(new_n627_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n671_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n491_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n547_), .B1(new_n494_), .B2(new_n501_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n629_), .A3(new_n662_), .ZN(new_n745_));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n700_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n742_), .A2(new_n747_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n740_), .B2(new_n490_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT48), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n749_), .A3(new_n490_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n740_), .B2(new_n689_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT49), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n745_), .A2(new_n754_), .A3(new_n689_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1334gat));
  AOI21_X1  g557(.A(new_n358_), .B1(new_n740_), .B2(new_n384_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n745_), .A2(new_n358_), .A3(new_n384_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n698_), .A2(new_n662_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n743_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n700_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n707_), .A2(new_n709_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n663_), .A2(new_n672_), .A3(new_n627_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n769_), .A2(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n700_), .A2(G85gat), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n767_), .A2(new_n768_), .B1(new_n773_), .B2(new_n774_), .ZN(G1336gat));
  AOI21_X1  g574(.A(G92gat), .B1(new_n765_), .B2(new_n490_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n490_), .A2(G92gat), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT116), .Z(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n773_), .B2(new_n778_), .ZN(G1337gat));
  XNOR2_X1  g578(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n689_), .B(new_n772_), .C1(new_n707_), .C2(new_n709_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(G99gat), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n781_), .A3(G99gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n765_), .A2(new_n499_), .A3(new_n568_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n780_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n785_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n787_), .B(new_n780_), .C1(new_n789_), .C2(new_n783_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n791_), .ZN(G1338gat));
  OAI211_X1 g591(.A(new_n384_), .B(new_n772_), .C1(new_n707_), .C2(new_n709_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(G106gat), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n743_), .A2(new_n384_), .A3(new_n569_), .A4(new_n764_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT119), .Z(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1339gat));
  AOI21_X1  g601(.A(new_n529_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n528_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n543_), .B1(new_n538_), .B2(new_n529_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n546_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n634_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n638_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n633_), .A2(new_n637_), .A3(KEYINPUT55), .A4(new_n634_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n645_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT56), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n645_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n808_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n808_), .B(KEYINPUT58), .C1(new_n814_), .C2(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n606_), .A3(new_n820_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n545_), .A2(new_n546_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n659_), .B2(new_n807_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n807_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT121), .B(new_n826_), .C1(new_n650_), .C2(new_n654_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n597_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n828_), .B2(new_n597_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n821_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n626_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n627_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n708_), .A2(new_n672_), .A3(new_n662_), .A4(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT54), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n700_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n547_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n819_), .A2(new_n606_), .A3(new_n820_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n828_), .A2(new_n597_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT57), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(new_n830_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT122), .B1(new_n848_), .B2(new_n835_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n833_), .A2(new_n850_), .A3(new_n627_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n851_), .A3(new_n837_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  INV_X1    g652(.A(new_n841_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n838_), .B2(new_n854_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n672_), .A3(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n844_), .B1(new_n857_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n662_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n842_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n855_), .A2(new_n662_), .A3(new_n856_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n859_), .ZN(G1341gat));
  NAND3_X1  g662(.A1(new_n842_), .A2(new_n207_), .A3(new_n835_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n855_), .A2(new_n626_), .A3(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n207_), .ZN(G1342gat));
  AOI21_X1  g665(.A(G134gat), .B1(new_n842_), .B2(new_n670_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n855_), .A2(new_n856_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT123), .B(G134gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n708_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n868_), .B2(new_n870_), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n288_), .A2(new_n384_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n491_), .A3(new_n490_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n838_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n547_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n663_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g677(.A1(new_n838_), .A2(new_n835_), .A3(new_n873_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(KEYINPUT124), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(KEYINPUT124), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n874_), .B2(new_n670_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n606_), .A2(G162gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT125), .Z(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n874_), .B2(new_n888_), .ZN(G1347gat));
  NAND2_X1  g688(.A1(new_n490_), .A2(new_n491_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n288_), .A2(new_n384_), .A3(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n852_), .A2(new_n547_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G169gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT126), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n895_), .A3(G169gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(KEYINPUT62), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n892_), .B2(G169gat), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  INV_X1    g698(.A(new_n892_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n899_), .B1(new_n900_), .B2(new_n234_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n901_), .ZN(G1348gat));
  NAND4_X1  g701(.A1(new_n838_), .A2(G176gat), .A3(new_n663_), .A4(new_n891_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT127), .Z(new_n904_));
  NAND2_X1  g703(.A1(new_n852_), .A2(new_n891_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n906_), .B2(new_n663_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n904_), .A2(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n905_), .A2(new_n244_), .A3(new_n626_), .ZN(new_n909_));
  INV_X1    g708(.A(G183gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n838_), .A2(new_n835_), .A3(new_n891_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n905_), .B2(new_n708_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n670_), .A2(new_n245_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n905_), .B2(new_n914_), .ZN(G1351gat));
  OR2_X1    g714(.A1(new_n872_), .A2(new_n890_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n839_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n547_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n663_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n338_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n326_), .B2(new_n920_), .ZN(G1353gat));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n625_), .A3(new_n623_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT63), .B(G211gat), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(new_n926_), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n917_), .A2(new_n928_), .A3(new_n670_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n839_), .A2(new_n708_), .A3(new_n916_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n928_), .ZN(G1355gat));
endmodule


