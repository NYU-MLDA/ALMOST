//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n988_, new_n989_, new_n991_,
    new_n992_, new_n994_, new_n996_, new_n997_, new_n998_, new_n1000_,
    new_n1001_, new_n1002_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT82), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT24), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT83), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(KEYINPUT84), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT84), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n216_), .B(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n221_), .B2(new_n214_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT24), .B1(new_n211_), .B2(new_n213_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n226_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n223_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT86), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n229_), .B2(KEYINPUT86), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT22), .B1(new_n209_), .B2(KEYINPUT85), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n209_), .A2(KEYINPUT22), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n210_), .B(new_n239_), .C1(new_n240_), .C2(KEYINPUT85), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n241_), .A2(new_n217_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n232_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT87), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT30), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n244_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT87), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n208_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n208_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G127gat), .B(G134gat), .Z(new_n254_));
  XOR2_X1   g053(.A(G113gat), .B(G120gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n253_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n251_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G1gat), .B(G29gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G85gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT0), .B(G57gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n256_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT3), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT2), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(KEYINPUT1), .B2(new_n276_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n276_), .A2(new_n279_), .A3(KEYINPUT1), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n276_), .B2(KEYINPUT1), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n278_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n270_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n272_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n269_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n282_), .A2(new_n284_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n256_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(KEYINPUT99), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT99), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n269_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT101), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT101), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n295_), .B(KEYINPUT100), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n286_), .A2(KEYINPUT4), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n268_), .B1(new_n302_), .B2(new_n308_), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n310_), .A2(new_n267_), .A3(new_n297_), .A4(new_n301_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT19), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G218gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G211gat), .ZN(new_n328_));
  INV_X1    g127(.A(G211gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G218gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n328_), .A2(new_n330_), .A3(new_n325_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n323_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n330_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT92), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(new_n325_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n321_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT21), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n335_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT21), .B1(new_n339_), .B2(new_n323_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT95), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n225_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n225_), .A2(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n224_), .A3(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT24), .A4(new_n216_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n235_), .A4(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT96), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n229_), .A2(new_n236_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G169gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n210_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n217_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT97), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n227_), .B(KEYINPUT23), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n237_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT97), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n217_), .A4(new_n354_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n350_), .A2(new_n351_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n235_), .A2(new_n349_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n362_), .A2(KEYINPUT96), .A3(new_n347_), .A4(new_n346_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n342_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT21), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(new_n340_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n244_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n320_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT98), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT98), .B(new_n320_), .C1(new_n364_), .C2(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n361_), .A2(new_n363_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(new_n367_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n244_), .A2(new_n367_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n320_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(KEYINPUT20), .A3(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n318_), .B1(new_n373_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n318_), .ZN(new_n382_));
  AOI211_X1 g181(.A(new_n382_), .B(new_n379_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n314_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n291_), .A2(KEYINPUT29), .ZN(new_n385_));
  INV_X1    g184(.A(G233gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n385_), .A2(new_n367_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n338_), .A2(new_n393_), .A3(new_n341_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT93), .B1(new_n366_), .B2(new_n340_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n394_), .A2(new_n395_), .B1(KEYINPUT29), .B2(new_n291_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n392_), .B1(new_n396_), .B2(new_n391_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n392_), .C1(new_n396_), .C2(new_n391_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT94), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n291_), .A2(KEYINPUT29), .ZN(new_n405_));
  XOR2_X1   g204(.A(G22gat), .B(G50gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT28), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n405_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n402_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n399_), .A2(new_n403_), .A3(new_n401_), .A4(new_n408_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n373_), .A2(new_n318_), .A3(new_n380_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n374_), .A2(new_n367_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n368_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(new_n320_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n358_), .A2(new_n217_), .A3(new_n354_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n394_), .A2(new_n395_), .A3(new_n350_), .A4(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT20), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT102), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT102), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT20), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n376_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n418_), .B1(new_n425_), .B2(new_n320_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n318_), .B(KEYINPUT103), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n414_), .B(KEYINPUT27), .C1(new_n426_), .C2(new_n427_), .ZN(new_n428_));
  AND4_X1   g227(.A1(new_n313_), .A2(new_n384_), .A3(new_n413_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n376_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n423_), .B1(new_n420_), .B2(KEYINPUT20), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n320_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n320_), .B2(new_n417_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n318_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n373_), .A2(new_n434_), .A3(new_n380_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n312_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n373_), .A2(new_n380_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n382_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n304_), .A2(new_n298_), .A3(new_n307_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n294_), .A2(new_n305_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n268_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT33), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n311_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n299_), .B(KEYINPUT101), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(KEYINPUT33), .A3(new_n267_), .A4(new_n310_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n440_), .A2(new_n445_), .A3(new_n414_), .A4(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n413_), .B1(new_n438_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n263_), .B1(new_n429_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n384_), .A2(new_n428_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n413_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n263_), .A2(new_n312_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G113gat), .B(G141gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT81), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G169gat), .B(G197gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT77), .B(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT14), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n462_), .B(new_n468_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n474_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(KEYINPUT15), .A3(new_n476_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n481_), .A2(new_n470_), .A3(new_n471_), .A4(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n479_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n477_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n470_), .A2(new_n486_), .A3(new_n471_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n479_), .B1(new_n478_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n461_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n484_), .A3(new_n460_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n456_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n495_));
  INV_X1    g294(.A(G71gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G78gat), .ZN(new_n497_));
  INV_X1    g296(.A(G78gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G71gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G57gat), .B(G64gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(KEYINPUT11), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n501_), .B2(KEYINPUT11), .ZN(new_n504_));
  INV_X1    g303(.A(G64gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G57gat), .ZN(new_n506_));
  INV_X1    g305(.A(G57gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G64gat), .ZN(new_n508_));
  AND4_X1   g307(.A1(new_n503_), .A2(new_n506_), .A3(new_n508_), .A4(KEYINPUT11), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n502_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n508_), .A3(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT68), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n506_), .A2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n506_), .A2(new_n508_), .A3(new_n503_), .A4(KEYINPUT11), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n512_), .A2(new_n515_), .A3(new_n500_), .A4(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n510_), .A2(new_n517_), .A3(KEYINPUT69), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT69), .B1(new_n510_), .B2(new_n517_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT6), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT67), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n529_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(new_n527_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n533_), .B1(new_n539_), .B2(new_n526_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT67), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n541_), .A3(KEYINPUT8), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT10), .B(G99gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n526_), .B1(new_n543_), .B2(G106gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545_));
  AND2_X1   g344(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n546_));
  NOR2_X1   g345(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(G92gat), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n531_), .A2(KEYINPUT9), .A3(new_n532_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(KEYINPUT66), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n552_), .A3(new_n549_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT67), .B1(new_n530_), .B2(new_n534_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT8), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n551_), .A2(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n521_), .A2(KEYINPUT70), .A3(new_n542_), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n510_), .A2(new_n517_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n518_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n535_), .A2(new_n536_), .A3(new_n555_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n550_), .A2(KEYINPUT66), .ZN(new_n564_));
  INV_X1    g363(.A(new_n544_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n553_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT8), .B1(new_n540_), .B2(KEYINPUT67), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n536_), .B(new_n533_), .C1(new_n539_), .C2(new_n526_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n563_), .B(new_n566_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n558_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n562_), .A2(new_n569_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n557_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT64), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n559_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n569_), .A2(new_n581_), .A3(KEYINPUT12), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n576_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n495_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n481_), .A2(new_n482_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n569_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n569_), .B2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT76), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n556_), .A2(new_n477_), .A3(new_n542_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT34), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT35), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT72), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n606_), .A2(KEYINPUT35), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n602_), .A2(new_n603_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n569_), .A2(new_n599_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT73), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n569_), .A2(new_n599_), .A3(new_n598_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n610_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT76), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n619_));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT75), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n608_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n609_), .B1(new_n569_), .B2(new_n486_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT74), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n626_), .B2(new_n602_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n618_), .A2(new_n619_), .A3(new_n623_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n619_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n623_), .A2(new_n619_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n603_), .B1(new_n602_), .B2(new_n610_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n615_), .A2(KEYINPUT76), .A3(new_n616_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT74), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n604_), .A2(new_n634_), .A3(new_n609_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n604_), .B2(new_n609_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n608_), .B1(new_n637_), .B2(new_n615_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n629_), .B(new_n630_), .C1(new_n633_), .C2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n628_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n628_), .A2(new_n639_), .A3(KEYINPUT37), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G127gat), .B(G155gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT17), .ZN(new_n650_));
  INV_X1    g449(.A(G231gat), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n386_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n470_), .A2(new_n471_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n521_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n562_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n650_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n649_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n656_), .A2(new_n581_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n559_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n659_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n644_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT80), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n494_), .A2(new_n597_), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n312_), .A3(new_n463_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n640_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n628_), .A2(new_n639_), .A3(KEYINPUT104), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n455_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n596_), .A2(new_n493_), .A3(new_n667_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n681_), .B2(new_n313_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n671_), .A2(new_n672_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n673_), .A2(new_n682_), .A3(new_n683_), .ZN(G1324gat));
  NAND3_X1  g483(.A1(new_n670_), .A2(new_n464_), .A3(new_n451_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(new_n451_), .A3(new_n680_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G8gat), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT39), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT39), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT40), .B(new_n685_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n681_), .B2(new_n263_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  INV_X1    g495(.A(new_n263_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n670_), .A2(new_n206_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n670_), .A2(new_n700_), .A3(new_n413_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n681_), .A2(new_n412_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n700_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(G1327gat));
  AND3_X1   g506(.A1(new_n628_), .A2(new_n639_), .A3(KEYINPUT104), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT104), .B1(new_n628_), .B2(new_n639_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n667_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n596_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n494_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n714_), .B2(new_n312_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n596_), .A2(new_n493_), .A3(new_n666_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n455_), .B2(new_n644_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n642_), .A2(new_n643_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT43), .B(new_n719_), .C1(new_n450_), .C2(new_n454_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n716_), .C1(new_n718_), .C2(new_n720_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n312_), .A2(G29gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n715_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n451_), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G36gat), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n451_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n384_), .A2(new_n428_), .A3(KEYINPUT106), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(G36gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n713_), .A2(KEYINPUT45), .A3(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT45), .B1(new_n713_), .B2(new_n736_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n729_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n729_), .A2(new_n739_), .A3(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1329gat));
  NAND4_X1  g543(.A1(new_n723_), .A2(G43gat), .A3(new_n697_), .A4(new_n724_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n203_), .B1(new_n713_), .B2(new_n263_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g547(.A1(new_n713_), .A2(G50gat), .A3(new_n412_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n725_), .B2(new_n413_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n723_), .A2(new_n750_), .A3(new_n413_), .A4(new_n724_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G50gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n751_), .B2(new_n753_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n456_), .A2(new_n492_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n596_), .A3(new_n669_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n507_), .B1(new_n756_), .B2(new_n313_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT108), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n493_), .A2(new_n666_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n597_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n678_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n507_), .A3(new_n313_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n758_), .A2(new_n764_), .ZN(G1332gat));
  INV_X1    g564(.A(new_n756_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n505_), .A3(new_n733_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n762_), .A2(new_n733_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(G64gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G64gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT110), .ZN(G1333gat));
  AOI21_X1  g572(.A(new_n496_), .B1(new_n762_), .B2(new_n697_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT49), .Z(new_n775_));
  NOR2_X1   g574(.A1(new_n263_), .A2(G71gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT111), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n756_), .B2(new_n777_), .ZN(G1334gat));
  AOI21_X1  g577(.A(new_n498_), .B1(new_n762_), .B2(new_n413_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT50), .Z(new_n780_));
  NAND3_X1  g579(.A1(new_n766_), .A2(new_n498_), .A3(new_n413_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n711_), .A2(new_n597_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n755_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT112), .B1(new_n755_), .B2(new_n783_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n312_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n718_), .A2(new_n720_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n597_), .A2(new_n492_), .A3(new_n666_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT113), .Z(new_n793_));
  NOR2_X1   g592(.A1(new_n546_), .A2(new_n547_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n313_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n789_), .B1(new_n793_), .B2(new_n795_), .ZN(G1336gat));
  AOI21_X1  g595(.A(G92gat), .B1(new_n788_), .B2(new_n451_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n733_), .A2(G92gat), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT114), .Z(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n793_), .B2(new_n799_), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n792_), .B2(new_n263_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n786_), .A2(new_n787_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n263_), .A2(new_n543_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n801_), .B(new_n805_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1338gat));
  NOR2_X1   g608(.A1(new_n412_), .A2(G106gat), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n413_), .B(new_n791_), .C1(new_n718_), .C2(new_n720_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(G106gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n812_), .B2(G106gat), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n802_), .A2(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  OAI221_X1 g617(.A(new_n818_), .B1(new_n814_), .B2(new_n815_), .C1(new_n802_), .C2(new_n811_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n594_), .A2(new_n590_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n478_), .A2(new_n487_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n479_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n478_), .A2(G229gat), .A3(new_n483_), .A4(G233gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n461_), .A3(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n491_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n590_), .A2(new_n492_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n557_), .A2(new_n570_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n542_), .A2(new_n556_), .B1(new_n561_), .B2(new_n518_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n582_), .B1(new_n832_), .B2(KEYINPUT12), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n575_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n578_), .A2(new_n580_), .A3(KEYINPUT55), .A4(new_n582_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n833_), .B2(new_n577_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n588_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n830_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n829_), .B1(new_n843_), .B2(KEYINPUT117), .ZN(new_n844_));
  INV_X1    g643(.A(new_n830_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n838_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n838_), .B2(new_n588_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT117), .B(new_n845_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n822_), .B1(new_n844_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n590_), .A2(new_n828_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT58), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n851_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(KEYINPUT118), .A3(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n644_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n850_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n848_), .A3(new_n829_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(new_n864_), .B2(new_n677_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n667_), .B1(new_n860_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT116), .B1(new_n493_), .B2(new_n666_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n869_));
  NOR4_X1   g668(.A1(new_n492_), .A2(new_n659_), .A3(new_n665_), .A4(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n871_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n867_), .B1(new_n719_), .B2(new_n872_), .ZN(new_n873_));
  AND4_X1   g672(.A1(new_n867_), .A2(new_n872_), .A3(new_n643_), .A4(new_n642_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n866_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n452_), .A2(new_n312_), .A3(new_n697_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G113gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n493_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n856_), .A2(KEYINPUT118), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n885_), .A2(KEYINPUT58), .B1(new_n643_), .B2(new_n642_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n886_), .A2(new_n858_), .B1(new_n864_), .B2(new_n822_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n677_), .B1(new_n844_), .B2(new_n849_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n821_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n666_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n884_), .B1(new_n890_), .B2(new_n875_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n866_), .A2(new_n876_), .A3(KEYINPUT119), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n879_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n881_), .B(new_n883_), .C1(new_n893_), .C2(new_n878_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT119), .B1(new_n866_), .B2(new_n876_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n492_), .B(new_n880_), .C1(new_n895_), .C2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n882_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n894_), .A2(new_n898_), .A3(KEYINPUT120), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1340gat));
  OAI21_X1  g702(.A(new_n881_), .B1(new_n893_), .B2(new_n878_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G120gat), .B1(new_n904_), .B2(new_n597_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n893_), .ZN(new_n906_));
  INV_X1    g705(.A(G120gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n597_), .B2(KEYINPUT60), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(KEYINPUT60), .B2(new_n907_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n905_), .B1(new_n906_), .B2(new_n909_), .ZN(G1341gat));
  OAI21_X1  g709(.A(G127gat), .B1(new_n904_), .B2(new_n667_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n667_), .A2(G127gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n906_), .B2(new_n912_), .ZN(G1342gat));
  OAI21_X1  g712(.A(G134gat), .B1(new_n904_), .B2(new_n719_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n677_), .A2(G134gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n906_), .B2(new_n915_), .ZN(G1343gat));
  AOI21_X1  g715(.A(new_n697_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n734_), .A2(new_n312_), .A3(new_n413_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  OR3_X1    g719(.A1(new_n920_), .A2(G141gat), .A3(new_n493_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G141gat), .B1(new_n920_), .B2(new_n493_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1344gat));
  INV_X1    g722(.A(new_n920_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT121), .B(G148gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n924_), .A2(new_n596_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n920_), .B2(new_n597_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1345gat));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G155gat), .ZN(new_n930_));
  OR3_X1    g729(.A1(new_n920_), .A2(new_n667_), .A3(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n920_), .B2(new_n667_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1346gat));
  NAND2_X1  g732(.A1(new_n644_), .A2(G162gat), .ZN(new_n934_));
  XOR2_X1   g733(.A(new_n934_), .B(KEYINPUT122), .Z(new_n935_));
  NAND3_X1  g734(.A1(new_n917_), .A2(new_n710_), .A3(new_n919_), .ZN(new_n936_));
  INV_X1    g735(.A(G162gat), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n924_), .A2(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(G1347gat));
  AND3_X1   g737(.A1(new_n384_), .A2(new_n428_), .A3(KEYINPUT106), .ZN(new_n939_));
  AOI21_X1  g738(.A(KEYINPUT106), .B1(new_n384_), .B2(new_n428_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n453_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  OAI211_X1 g742(.A(KEYINPUT123), .B(new_n453_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n877_), .A2(new_n412_), .A3(new_n945_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n946_), .A2(KEYINPUT127), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(KEYINPUT127), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n947_), .A2(new_n353_), .A3(new_n492_), .A4(new_n948_), .ZN(new_n949_));
  AOI211_X1 g748(.A(new_n413_), .B(new_n493_), .C1(new_n943_), .C2(new_n944_), .ZN(new_n950_));
  AOI21_X1  g749(.A(KEYINPUT124), .B1(new_n877_), .B2(new_n950_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n861_), .A2(new_n862_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n710_), .B1(new_n952_), .B2(new_n848_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n850_), .B(new_n859_), .C1(new_n953_), .C2(KEYINPUT57), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n875_), .B1(new_n954_), .B2(new_n667_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956_));
  AOI21_X1  g755(.A(KEYINPUT123), .B1(new_n733_), .B2(new_n453_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n944_), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n412_), .B(new_n492_), .C1(new_n957_), .C2(new_n958_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n955_), .A2(new_n956_), .A3(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G169gat), .B1(new_n951_), .B2(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n961_), .A2(new_n962_), .A3(KEYINPUT62), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n956_), .B1(new_n955_), .B2(new_n959_), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n950_), .B(KEYINPUT124), .C1(new_n890_), .C2(new_n875_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n209_), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967_));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n963_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n964_), .A2(new_n965_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n209_), .A2(KEYINPUT62), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n970_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n972_), .ZN(new_n974_));
  AOI211_X1 g773(.A(KEYINPUT125), .B(new_n974_), .C1(new_n964_), .C2(new_n965_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n973_), .A2(new_n975_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n949_), .B1(new_n969_), .B2(new_n976_), .ZN(G1348gat));
  NAND3_X1  g776(.A1(new_n947_), .A2(new_n596_), .A3(new_n948_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n413_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n979_));
  AOI211_X1 g778(.A(new_n210_), .B(new_n597_), .C1(new_n943_), .C2(new_n944_), .ZN(new_n980_));
  AOI22_X1  g779(.A1(new_n978_), .A2(new_n210_), .B1(new_n979_), .B2(new_n980_), .ZN(G1349gat));
  NAND2_X1  g780(.A1(new_n947_), .A2(new_n948_), .ZN(new_n982_));
  INV_X1    g781(.A(new_n982_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n667_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n984_));
  INV_X1    g783(.A(G183gat), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n979_), .A2(new_n666_), .A3(new_n945_), .ZN(new_n986_));
  AOI22_X1  g785(.A1(new_n983_), .A2(new_n984_), .B1(new_n985_), .B2(new_n986_), .ZN(G1350gat));
  OAI21_X1  g786(.A(G190gat), .B1(new_n982_), .B2(new_n719_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n710_), .A2(new_n224_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n988_), .B1(new_n982_), .B2(new_n989_), .ZN(G1351gat));
  NOR3_X1   g789(.A1(new_n734_), .A2(new_n312_), .A3(new_n412_), .ZN(new_n991_));
  NAND3_X1  g790(.A1(new_n917_), .A2(new_n492_), .A3(new_n991_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g792(.A1(new_n917_), .A2(new_n596_), .A3(new_n991_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n994_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g794(.A(KEYINPUT63), .B(G211gat), .ZN(new_n996_));
  OR2_X1    g795(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n997_));
  NAND3_X1  g796(.A1(new_n917_), .A2(new_n666_), .A3(new_n991_), .ZN(new_n998_));
  MUX2_X1   g797(.A(new_n996_), .B(new_n997_), .S(new_n998_), .Z(G1354gat));
  NAND2_X1  g798(.A1(new_n917_), .A2(new_n991_), .ZN(new_n1000_));
  OAI21_X1  g799(.A(G218gat), .B1(new_n1000_), .B2(new_n719_), .ZN(new_n1001_));
  NAND2_X1  g800(.A1(new_n710_), .A2(new_n327_), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n1000_), .B2(new_n1002_), .ZN(G1355gat));
endmodule


