//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n974_, new_n975_, new_n976_, new_n978_,
    new_n979_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n989_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n1000_,
    new_n1001_, new_n1002_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(KEYINPUT1), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n209_), .A3(KEYINPUT1), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n208_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n206_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n210_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(new_n213_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT87), .B1(new_n216_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n212_), .A2(new_n213_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n211_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n215_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n207_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT87), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n223_), .A2(new_n225_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235_));
  XOR2_X1   g034(.A(G127gat), .B(G134gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n227_), .A2(new_n234_), .A3(new_n235_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n227_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n231_), .A2(new_n233_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(new_n238_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT4), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n244_), .A2(new_n246_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n243_), .A2(new_n247_), .B1(new_n248_), .B2(new_n240_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G57gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT95), .B1(new_n249_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT94), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n249_), .A2(new_n255_), .A3(new_n253_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(new_n241_), .A3(new_n239_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n244_), .A2(new_n246_), .A3(new_n240_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT95), .ZN(new_n260_));
  INV_X1    g059(.A(new_n253_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT4), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n258_), .B(new_n253_), .C1(new_n263_), .C2(new_n242_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT94), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n254_), .A2(new_n256_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(G197gat), .A2(G204gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT88), .B1(new_n273_), .B2(KEYINPUT21), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n275_), .B(new_n269_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n270_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT89), .ZN(new_n278_));
  INV_X1    g077(.A(G218gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G211gat), .ZN(new_n280_));
  INV_X1    g079(.A(G211gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G218gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n273_), .B2(KEYINPUT21), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n275_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n276_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n268_), .A2(new_n269_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n283_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n278_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT22), .B(G169gat), .ZN(new_n293_));
  INV_X1    g092(.A(G176gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n296_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(G169gat), .B2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(G169gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n294_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n309_), .A3(new_n294_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n303_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT91), .B1(new_n292_), .B2(new_n315_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n287_), .A2(new_n288_), .B1(new_n290_), .B2(new_n283_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT91), .ZN(new_n318_));
  INV_X1    g117(.A(new_n315_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n278_), .A4(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT20), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT22), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G169gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(G176gat), .B1(new_n326_), .B2(KEYINPUT82), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(KEYINPUT82), .B2(new_n293_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n327_), .B(KEYINPUT83), .C1(KEYINPUT82), .C2(new_n293_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n302_), .A2(new_n296_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n312_), .A2(KEYINPUT81), .ZN(new_n334_));
  INV_X1    g133(.A(new_n314_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n304_), .A2(new_n305_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n333_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n339_));
  AOI211_X1 g138(.A(new_n322_), .B(new_n324_), .C1(new_n292_), .C2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n314_), .B1(new_n312_), .B2(KEYINPUT81), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(KEYINPUT81), .B2(new_n312_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(new_n317_), .A3(new_n333_), .A4(new_n278_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n291_), .B1(new_n277_), .B2(KEYINPUT89), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n287_), .A2(new_n288_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n315_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(KEYINPUT20), .A3(new_n346_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n321_), .A2(new_n340_), .B1(new_n347_), .B2(new_n324_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n324_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n343_), .A2(new_n346_), .A3(KEYINPUT20), .A4(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n322_), .B1(new_n292_), .B2(new_n339_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n315_), .A2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n303_), .B(KEYINPUT93), .C1(new_n312_), .C2(new_n314_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n317_), .A2(new_n361_), .A3(new_n278_), .A4(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n356_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT32), .B(new_n353_), .C1(new_n358_), .C2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n266_), .A2(new_n355_), .A3(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n264_), .B(KEYINPUT33), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n321_), .A2(new_n340_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n347_), .A2(new_n324_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n353_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n352_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n244_), .A2(new_n246_), .A3(new_n241_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n261_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(KEYINPUT92), .A3(new_n261_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n247_), .A2(new_n240_), .A3(new_n239_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n367_), .A2(new_n370_), .A3(new_n372_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n366_), .A2(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n317_), .A2(new_n278_), .B1(KEYINPUT29), .B2(new_n245_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT90), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n245_), .A2(KEYINPUT29), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n292_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n387_));
  INV_X1    g186(.A(new_n383_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n227_), .A2(new_n234_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n383_), .B(new_n292_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G78gat), .B(G106gat), .Z(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT28), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n397_), .A2(KEYINPUT28), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G22gat), .B(G50gat), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n395_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n390_), .A2(new_n405_), .A3(new_n393_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n396_), .A2(new_n403_), .A3(new_n404_), .A4(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n390_), .A2(new_n405_), .A3(new_n393_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n401_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n400_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n398_), .ZN(new_n412_));
  OAI22_X1  g211(.A1(new_n408_), .A2(new_n409_), .B1(new_n402_), .B2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n266_), .B1(new_n407_), .B2(new_n413_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT96), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n352_), .C1(new_n358_), .C2(new_n364_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n370_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n292_), .A2(new_n339_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n363_), .A3(KEYINPUT20), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n324_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n357_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n416_), .B1(new_n422_), .B2(new_n352_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT27), .B1(new_n418_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n372_), .A2(new_n425_), .A3(new_n370_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n381_), .A2(new_n414_), .B1(new_n415_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n339_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G43gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(G15gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n436_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n430_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n443_), .B2(KEYINPUT85), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n440_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n444_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n202_), .B1(new_n428_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n355_), .A2(new_n365_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n253_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n454_), .A2(new_n260_), .B1(new_n264_), .B2(KEYINPUT94), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n454_), .A2(new_n260_), .B1(new_n264_), .B2(KEYINPUT94), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n453_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n372_), .A2(new_n370_), .A3(new_n379_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n264_), .B(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n414_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n415_), .A2(new_n427_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n447_), .A2(new_n450_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT97), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n407_), .A2(new_n413_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n266_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n427_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n452_), .A2(new_n467_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  INV_X1    g272(.A(G1gat), .ZN(new_n474_));
  INV_X1    g273(.A(G8gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G29gat), .B(G36gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n479_), .B(new_n482_), .Z(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n482_), .B(KEYINPUT15), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n479_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n479_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(new_n482_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n483_), .A2(new_n485_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G113gat), .B(G141gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT79), .ZN(new_n492_));
  XOR2_X1   g291(.A(G169gat), .B(G197gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n490_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT80), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n472_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G190gat), .B(G218gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G134gat), .B(G162gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT36), .Z(new_n501_));
  INV_X1    g300(.A(G85gat), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT64), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT64), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT9), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n504_), .A2(new_n506_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n505_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n510_), .A2(new_n513_), .A3(new_n517_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT65), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n518_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n517_), .A4(new_n510_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n520_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529_));
  INV_X1    g328(.A(G99gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n515_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n523_), .A3(new_n524_), .A4(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  INV_X1    g333(.A(new_n509_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n534_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT69), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n538_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT8), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT69), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n528_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n486_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n520_), .B(new_n527_), .C1(new_n540_), .C2(new_n539_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT75), .B1(new_n550_), .B2(new_n482_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(new_n552_), .B2(KEYINPUT74), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n548_), .A2(new_n551_), .A3(new_n560_), .A4(new_n557_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n556_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n554_), .A3(new_n561_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n501_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n555_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n500_), .A2(KEYINPUT36), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n563_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n565_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n501_), .B(KEYINPUT76), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n570_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT77), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n569_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n572_), .B1(new_n567_), .B2(new_n563_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT37), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n565_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G71gat), .B(G78gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT67), .ZN(new_n585_));
  INV_X1    g384(.A(G57gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(G64gat), .ZN(new_n587_));
  INV_X1    g386(.A(G64gat), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(G57gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(G57gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(G64gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT67), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n584_), .B1(new_n594_), .B2(KEYINPUT11), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n594_), .B2(KEYINPUT11), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT11), .ZN(new_n598_));
  AOI211_X1 g397(.A(KEYINPUT68), .B(new_n598_), .C1(new_n590_), .C2(new_n593_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT67), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT67), .B1(new_n591_), .B2(new_n592_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n583_), .B1(new_n603_), .B2(new_n598_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT11), .B1(new_n601_), .B2(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT68), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n594_), .A2(new_n596_), .A3(KEYINPUT11), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n549_), .B1(new_n600_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n600_), .A2(new_n549_), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n608_), .A4(new_n600_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n616_), .A2(new_n613_), .A3(new_n610_), .A4(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(G176gat), .B(G204gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT71), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT72), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n621_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n619_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT13), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT13), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n479_), .B(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n600_), .A2(new_n608_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT17), .ZN(new_n639_));
  XOR2_X1   g438(.A(G127gat), .B(G155gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n638_), .A2(new_n639_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(KEYINPUT17), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n638_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n576_), .A2(new_n582_), .A3(new_n634_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n497_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n266_), .A2(KEYINPUT98), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n266_), .A2(KEYINPUT98), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(new_n474_), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n565_), .A2(new_n569_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n451_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n471_), .B1(new_n661_), .B2(KEYINPUT97), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n428_), .A2(new_n202_), .A3(new_n451_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT99), .B(new_n660_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT99), .B1(new_n472_), .B2(new_n660_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n495_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n633_), .A2(new_n668_), .A3(new_n648_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n266_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G1gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n659_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1324gat));
  INV_X1    g474(.A(new_n427_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n653_), .A2(new_n475_), .A3(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n676_), .B(new_n669_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(G8gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n678_), .B2(G8gat), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT39), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n678_), .A2(G8gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT101), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(new_n680_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n677_), .B1(new_n683_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n677_), .B(new_n689_), .C1(new_n683_), .C2(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1325gat));
  NAND3_X1  g492(.A1(new_n653_), .A2(new_n438_), .A3(new_n451_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n667_), .A2(new_n451_), .A3(new_n669_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n695_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n695_), .B2(G15gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n653_), .A2(new_n700_), .A3(new_n468_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n670_), .A2(new_n468_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G22gat), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT42), .B(new_n700_), .C1(new_n670_), .C2(new_n468_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1327gat));
  NOR3_X1   g505(.A1(new_n633_), .A2(new_n660_), .A3(new_n649_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n497_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n266_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n633_), .A2(new_n668_), .A3(new_n649_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n576_), .A2(new_n582_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n712_), .B(new_n713_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n712_), .B1(new_n472_), .B2(new_n713_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n711_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n711_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n713_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT43), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n714_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(G29gat), .A3(new_n657_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n723_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n711_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730_));
  INV_X1    g529(.A(new_n727_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n729_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n710_), .B1(new_n726_), .B2(new_n733_), .ZN(G1328gat));
  XNOR2_X1  g533(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n717_), .A2(new_n718_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n676_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n728_), .A2(new_n732_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G36gat), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n708_), .A2(G36gat), .A3(new_n427_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT45), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n735_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(G36gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n427_), .B1(new_n719_), .B2(new_n724_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n733_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n735_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n747_), .A2(new_n742_), .A3(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n744_), .A2(new_n749_), .ZN(G1329gat));
  NAND4_X1  g549(.A1(new_n733_), .A2(new_n725_), .A3(G43gat), .A4(new_n451_), .ZN(new_n751_));
  INV_X1    g550(.A(G43gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n708_), .B2(new_n466_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1330gat));
  AOI21_X1  g556(.A(G50gat), .B1(new_n709_), .B2(new_n468_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n725_), .A2(G50gat), .A3(new_n468_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n733_), .ZN(G1331gat));
  NOR3_X1   g559(.A1(new_n634_), .A2(new_n648_), .A3(new_n496_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n667_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G57gat), .B1(new_n763_), .B2(new_n470_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n472_), .A2(new_n668_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n634_), .B1(new_n765_), .B2(KEYINPUT109), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n472_), .A2(new_n767_), .A3(new_n668_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n713_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n649_), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n586_), .A3(new_n657_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(new_n772_), .ZN(G1332gat));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n588_), .A3(new_n676_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n762_), .A2(new_n676_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G64gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT48), .B(new_n588_), .C1(new_n762_), .C2(new_n676_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n771_), .A2(new_n780_), .A3(new_n451_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n762_), .A2(new_n451_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G71gat), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT49), .B(new_n780_), .C1(new_n762_), .C2(new_n451_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n771_), .A2(new_n787_), .A3(new_n468_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n762_), .A2(new_n468_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(G78gat), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G78gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n660_), .A2(new_n649_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n769_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n502_), .A3(new_n657_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n722_), .A2(new_n714_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n634_), .A2(new_n495_), .A3(new_n649_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n799_), .A2(KEYINPUT111), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(KEYINPUT111), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n470_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n796_), .B1(new_n804_), .B2(new_n502_), .ZN(G1336gat));
  NAND3_X1  g604(.A1(new_n795_), .A2(new_n503_), .A3(new_n676_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n427_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n503_), .ZN(G1337gat));
  AND3_X1   g607(.A1(new_n451_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n769_), .A2(new_n794_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT51), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n451_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G99gat), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n811_), .A2(KEYINPUT51), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n816_), .B(new_n813_), .C1(new_n814_), .C2(G99gat), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1338gat));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n797_), .A2(new_n468_), .A3(new_n798_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(G106gat), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(G106gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(KEYINPUT114), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n824_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n414_), .A2(G106gat), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n766_), .A2(new_n794_), .A3(new_n768_), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .A4(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n826_), .A2(KEYINPUT114), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n835_), .A2(new_n824_), .A3(new_n823_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n829_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n838_), .ZN(G1339gat));
  NAND3_X1  g638(.A1(new_n657_), .A2(new_n427_), .A3(new_n469_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n660_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n494_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n484_), .B1(new_n488_), .B2(new_n482_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n487_), .A2(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n490_), .A2(new_n494_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n495_), .A2(new_n627_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT115), .B1(new_n619_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n619_), .A2(new_n850_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n609_), .B1(new_n617_), .B2(new_n611_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n616_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n614_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n619_), .A2(KEYINPUT115), .A3(new_n850_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n626_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n613_), .B1(new_n853_), .B2(new_n616_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n850_), .B2(new_n619_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n616_), .A2(new_n610_), .A3(new_n618_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(KEYINPUT55), .A4(new_n613_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n861_), .A2(new_n862_), .A3(new_n865_), .A4(new_n851_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n858_), .A2(new_n859_), .A3(new_n866_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n865_), .A2(new_n851_), .A3(new_n852_), .A4(new_n855_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n626_), .B1(new_n871_), .B2(KEYINPUT116), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT56), .A3(new_n866_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n849_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n848_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n849_), .ZN(new_n877_));
  AND4_X1   g676(.A1(KEYINPUT56), .A2(new_n858_), .A3(new_n859_), .A4(new_n866_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n868_), .B1(new_n872_), .B2(new_n866_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n875_), .B(new_n877_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n843_), .B1(new_n876_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n627_), .A2(new_n847_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n867_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n873_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT58), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n886_), .A2(KEYINPUT58), .B1(new_n576_), .B2(new_n582_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n882_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT118), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n880_), .A3(new_n848_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n893_), .B2(new_n660_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n648_), .B1(new_n890_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n896_));
  INV_X1    g695(.A(new_n496_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n651_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT54), .B1(new_n650_), .B2(new_n496_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n840_), .B1(new_n895_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n495_), .ZN(new_n902_));
  INV_X1    g701(.A(G113gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT119), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n906_), .A3(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT120), .B1(new_n901_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n898_), .A2(new_n899_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n660_), .B1(new_n876_), .B2(new_n881_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n842_), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n893_), .A2(new_n843_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n912_), .B1(new_n916_), .B2(new_n648_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n911_), .B(KEYINPUT59), .C1(new_n917_), .C2(new_n840_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n840_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n649_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n909_), .B(new_n920_), .C1(new_n921_), .C2(new_n912_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n895_), .A2(new_n900_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n925_), .A2(KEYINPUT121), .A3(new_n909_), .A4(new_n920_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n919_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n897_), .A2(new_n903_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n908_), .B1(new_n928_), .B2(new_n929_), .ZN(G1340gat));
  NAND3_X1  g729(.A1(new_n919_), .A2(new_n927_), .A3(new_n633_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G120gat), .ZN(new_n932_));
  INV_X1    g731(.A(G120gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n634_), .B2(KEYINPUT60), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n901_), .B(new_n934_), .C1(KEYINPUT60), .C2(new_n933_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n935_), .ZN(G1341gat));
  NAND3_X1  g735(.A1(new_n919_), .A2(new_n927_), .A3(new_n649_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G127gat), .ZN(new_n938_));
  INV_X1    g737(.A(G127gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n901_), .A2(new_n939_), .A3(new_n649_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1342gat));
  AOI21_X1  g740(.A(G134gat), .B1(new_n901_), .B2(new_n841_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT122), .B(G134gat), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n770_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n942_), .B1(new_n928_), .B2(new_n944_), .ZN(G1343gat));
  NOR3_X1   g744(.A1(new_n676_), .A2(new_n451_), .A3(new_n414_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n925_), .A2(new_n657_), .A3(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n668_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n203_), .ZN(G1344gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n634_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT123), .B(G148gat), .Z(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1345gat));
  NOR2_X1   g751(.A1(new_n947_), .A2(new_n648_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT61), .B(G155gat), .Z(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1346gat));
  OAI21_X1  g754(.A(G162gat), .B1(new_n947_), .B2(new_n770_), .ZN(new_n956_));
  OR2_X1    g755(.A1(new_n660_), .A2(G162gat), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n947_), .B2(new_n957_), .ZN(G1347gat));
  NOR3_X1   g757(.A1(new_n657_), .A2(new_n466_), .A3(new_n427_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n925_), .A2(new_n414_), .A3(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G169gat), .B1(new_n960_), .B2(new_n668_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962_));
  OR2_X1    g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n960_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n964_), .A2(new_n293_), .A3(new_n495_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n961_), .A2(new_n962_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n963_), .A2(new_n965_), .A3(new_n966_), .ZN(G1348gat));
  AOI21_X1  g766(.A(G176gat), .B1(new_n964_), .B2(new_n633_), .ZN(new_n968_));
  OR3_X1    g767(.A1(new_n917_), .A2(KEYINPUT124), .A3(new_n468_), .ZN(new_n969_));
  OAI21_X1  g768(.A(KEYINPUT124), .B1(new_n917_), .B2(new_n468_), .ZN(new_n970_));
  AND2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  AND3_X1   g770(.A1(new_n959_), .A2(G176gat), .A3(new_n633_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n968_), .B1(new_n971_), .B2(new_n972_), .ZN(G1349gat));
  NOR3_X1   g772(.A1(new_n960_), .A2(new_n304_), .A3(new_n648_), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n969_), .A2(new_n649_), .A3(new_n959_), .A4(new_n970_), .ZN(new_n975_));
  INV_X1    g774(.A(G183gat), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n974_), .B1(new_n975_), .B2(new_n976_), .ZN(G1350gat));
  OAI21_X1  g776(.A(G190gat), .B1(new_n960_), .B2(new_n770_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n841_), .A2(new_n305_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n960_), .B2(new_n979_), .ZN(G1351gat));
  NAND3_X1  g779(.A1(new_n676_), .A2(new_n466_), .A3(new_n415_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n917_), .A2(new_n981_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n495_), .ZN(new_n983_));
  INV_X1    g782(.A(G197gat), .ZN(new_n984_));
  AND3_X1   g783(.A1(new_n983_), .A2(KEYINPUT125), .A3(new_n984_), .ZN(new_n985_));
  AOI21_X1  g784(.A(KEYINPUT125), .B1(new_n983_), .B2(new_n984_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n983_), .A2(new_n984_), .ZN(new_n987_));
  NOR3_X1   g786(.A1(new_n985_), .A2(new_n986_), .A3(new_n987_), .ZN(G1352gat));
  NAND2_X1  g787(.A1(new_n982_), .A2(new_n633_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(new_n989_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g789(.A1(new_n982_), .A2(new_n649_), .ZN(new_n991_));
  XNOR2_X1  g790(.A(KEYINPUT63), .B(G211gat), .ZN(new_n992_));
  NOR2_X1   g791(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n991_), .A2(new_n994_), .A3(new_n281_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n995_), .A2(KEYINPUT126), .ZN(new_n996_));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n997_));
  NAND4_X1  g796(.A1(new_n991_), .A2(new_n997_), .A3(new_n994_), .A4(new_n281_), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n993_), .B1(new_n996_), .B2(new_n998_), .ZN(G1354gat));
  AOI21_X1  g798(.A(G218gat), .B1(new_n982_), .B2(new_n841_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n713_), .A2(G218gat), .ZN(new_n1001_));
  XNOR2_X1  g800(.A(new_n1001_), .B(KEYINPUT127), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n1000_), .B1(new_n982_), .B2(new_n1002_), .ZN(G1355gat));
endmodule


