//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n205_), .A2(new_n209_), .B1(new_n212_), .B2(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n215_), .A2(new_n217_), .B1(new_n210_), .B2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n213_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n221_));
  INV_X1    g020(.A(new_n208_), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n206_), .ZN(new_n225_));
  AND4_X1   g024(.A1(KEYINPUT65), .A2(new_n221_), .A3(new_n219_), .A4(new_n225_), .ZN(new_n226_));
  OAI22_X1  g025(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n216_), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n227_), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G85gat), .B(G92gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(KEYINPUT67), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n220_), .A2(new_n226_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(new_n225_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n219_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n213_), .A2(KEYINPUT65), .A3(new_n219_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n233_), .A2(new_n236_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n251_), .A3(KEYINPUT68), .ZN(new_n252_));
  INV_X1    g051(.A(G64gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G57gat), .ZN(new_n254_));
  INV_X1    g053(.A(G57gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G64gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT69), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n254_), .B2(new_n256_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT11), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n255_), .A2(G64gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n253_), .A2(G57gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT69), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G71gat), .B(G78gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT11), .B(new_n267_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT70), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n241_), .A2(new_n252_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n275_), .A2(KEYINPUT71), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n241_), .A2(new_n252_), .A3(new_n272_), .A4(new_n274_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n275_), .B2(KEYINPUT71), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n204_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT72), .B1(new_n275_), .B2(KEYINPUT12), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n272_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n239_), .A2(new_n240_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT68), .B1(new_n247_), .B2(new_n251_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n273_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n239_), .A3(KEYINPUT12), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n282_), .A2(new_n283_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n281_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n280_), .A2(new_n287_), .A3(new_n293_), .A4(new_n203_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n279_), .A2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G120gat), .B(G148gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G176gat), .B(G204gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n279_), .A2(new_n294_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n301_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n295_), .A2(new_n302_), .A3(new_n300_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n202_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT13), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G29gat), .B(G36gat), .Z(new_n313_));
  XOR2_X1   g112(.A(G43gat), .B(G50gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(G1gat), .A2(G8gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G1gat), .A2(G8gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT78), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G15gat), .ZN(new_n323_));
  INV_X1    g122(.A(G22gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G15gat), .A2(G22gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT14), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n325_), .A2(new_n326_), .B1(new_n327_), .B2(new_n317_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n320_), .B(KEYINPUT79), .ZN(new_n330_));
  INV_X1    g129(.A(new_n328_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n316_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n331_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n322_), .A2(new_n328_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n315_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(KEYINPUT82), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n335_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n316_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n315_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n338_), .A3(new_n336_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n346_), .A2(KEYINPUT83), .A3(new_n338_), .A4(new_n336_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n343_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G113gat), .B(G141gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT84), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G169gat), .B(G197gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n343_), .A2(new_n349_), .A3(new_n350_), .A4(new_n355_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n312_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT88), .B(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G71gat), .B(G99gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT86), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT25), .B(G183gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT26), .B(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n369_), .A2(new_n372_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT24), .ZN(new_n379_));
  OAI221_X1 g178(.A(new_n377_), .B1(new_n376_), .B2(new_n375_), .C1(new_n372_), .C2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(G183gat), .B2(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT87), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n384_), .B2(new_n381_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G169gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n384_), .B2(KEYINPUT23), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n386_), .A2(KEYINPUT30), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT30), .B1(new_n386_), .B2(new_n393_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n368_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n386_), .A2(new_n393_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(KEYINPUT89), .A3(new_n394_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n367_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT89), .B1(new_n400_), .B2(new_n394_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n367_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G127gat), .B(G134gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT31), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n402_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n395_), .A2(new_n396_), .A3(new_n368_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n404_), .B1(new_n412_), .B2(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n397_), .A2(new_n367_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G155gat), .B(G162gat), .Z(new_n417_));
  OR2_X1    g216(.A1(G141gat), .A2(G148gat), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n418_), .A2(KEYINPUT3), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G141gat), .A2(G148gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT2), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(KEYINPUT3), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT90), .Z(new_n426_));
  OAI21_X1  g225(.A(new_n417_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT1), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n417_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n420_), .A4(new_n418_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n432_), .A2(KEYINPUT29), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT28), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G22gat), .B(G50gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(KEYINPUT28), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n437_), .A2(new_n440_), .A3(KEYINPUT91), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT92), .B(G197gat), .Z(new_n446_));
  INV_X1    g245(.A(G204gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT21), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(G197gat), .B2(G204gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(G204gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT93), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(G197gat), .B2(new_n447_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n451_), .B(new_n452_), .C1(new_n457_), .C2(KEYINPUT21), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n449_), .B1(new_n452_), .B2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n457_), .B(new_n460_), .C1(new_n459_), .C2(new_n452_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n432_), .A2(KEYINPUT29), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT95), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G78gat), .B(G106gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT96), .Z(new_n469_));
  OAI211_X1 g268(.A(new_n462_), .B(new_n463_), .C1(KEYINPUT95), .C2(new_n465_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n467_), .A2(KEYINPUT97), .A3(new_n470_), .A4(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n467_), .A2(new_n470_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n445_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n477_), .A2(new_n471_), .A3(new_n437_), .A4(new_n440_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n416_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n479_), .B(new_n480_), .C1(new_n411_), .C2(new_n415_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n432_), .B(new_n408_), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT4), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G225gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n432_), .A2(new_n408_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n486_), .B(new_n488_), .C1(KEYINPUT4), .C2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G85gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT0), .B(G57gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n487_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT101), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT101), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n485_), .A2(new_n497_), .A3(new_n487_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n490_), .A2(new_n494_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT103), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n496_), .A2(new_n498_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT103), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n494_), .A4(new_n490_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n490_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n494_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT104), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT22), .B(G169gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT100), .ZN(new_n510_));
  OAI221_X1 g309(.A(new_n378_), .B1(new_n385_), .B2(new_n392_), .C1(G176gat), .C2(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n378_), .A2(KEYINPUT99), .A3(KEYINPUT24), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT99), .B1(new_n378_), .B2(KEYINPUT24), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n372_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n370_), .A2(new_n369_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n390_), .A2(new_n375_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n511_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n462_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(KEYINPUT20), .C1(new_n398_), .C2(new_n462_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G226gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G8gat), .B(G36gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT18), .ZN(new_n525_));
  XOR2_X1   g324(.A(G64gat), .B(G92gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n398_), .A2(new_n462_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n462_), .A2(new_n517_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n522_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT20), .A4(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT105), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n523_), .A2(new_n531_), .A3(KEYINPUT105), .A4(new_n527_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n462_), .B2(new_n517_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n386_), .A2(new_n393_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n522_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n538_), .B(KEYINPUT102), .C1(new_n522_), .C2(new_n519_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT102), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n540_), .B(new_n522_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n534_), .B(new_n535_), .C1(new_n542_), .C2(new_n527_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT27), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n523_), .A2(new_n531_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n527_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT27), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n484_), .A2(new_n508_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n481_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n501_), .A2(KEYINPUT33), .A3(new_n494_), .A4(new_n490_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n486_), .B1(KEYINPUT4), .B2(new_n489_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(new_n488_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n485_), .A2(new_n488_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n505_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT33), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n499_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n546_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n507_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n527_), .A2(KEYINPUT32), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n523_), .A2(new_n531_), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n542_), .B2(new_n561_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n416_), .B(new_n551_), .C1(new_n559_), .C2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n550_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n361_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT36), .Z(new_n571_));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT34), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n345_), .A2(new_n239_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n241_), .A2(new_n252_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n316_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n572_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n571_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n570_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT77), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT80), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n340_), .B(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(new_n292_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n292_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT16), .ZN(new_n602_));
  XOR2_X1   g401(.A(G183gat), .B(G211gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT17), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n600_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n598_), .B(KEYINPUT81), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n288_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n604_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n607_), .B2(new_n273_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n606_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n595_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT106), .B1(new_n567_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT106), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n361_), .A2(new_n617_), .A3(new_n566_), .A4(new_n614_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n508_), .A2(G1gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n616_), .A2(KEYINPUT38), .A3(new_n618_), .A4(new_n619_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n587_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n613_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n567_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n508_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G1gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(new_n623_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(G8gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n549_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n616_), .A2(new_n634_), .A3(new_n635_), .A4(new_n618_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n627_), .A2(new_n635_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(G8gat), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT39), .B(new_n634_), .C1(new_n627_), .C2(new_n635_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n641_), .B(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(new_n416_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n323_), .B1(new_n627_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n616_), .A2(new_n618_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n323_), .A3(new_n645_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n647_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(G1326gat));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n324_), .A3(new_n481_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n627_), .A2(new_n481_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G22gat), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT42), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT42), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(new_n613_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n567_), .A2(new_n659_), .A3(new_n587_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n628_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT110), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT44), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n595_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n550_), .B2(new_n565_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n595_), .A2(KEYINPUT109), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n595_), .A2(KEYINPUT109), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n566_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n667_), .B1(new_n671_), .B2(KEYINPUT43), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n361_), .A2(new_n613_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n664_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n666_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n566_), .A2(new_n675_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n550_), .A2(new_n565_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n665_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n673_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n663_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n628_), .A2(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n661_), .B1(new_n681_), .B2(new_n682_), .ZN(G1328gat));
  NAND2_X1  g482(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n672_), .A2(new_n664_), .A3(new_n673_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n663_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n635_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G36gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n659_), .A2(new_n587_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n549_), .A2(G36gat), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n361_), .A2(new_n566_), .A3(new_n690_), .A4(new_n691_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT45), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(KEYINPUT45), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n689_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n684_), .B1(new_n688_), .B2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n549_), .B1(new_n674_), .B2(new_n680_), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n684_), .B(new_n695_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(G1329gat));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n645_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G43gat), .ZN(new_n704_));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n660_), .A2(new_n705_), .A3(new_n645_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n416_), .B1(new_n674_), .B2(new_n680_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n702_), .B(new_n706_), .C1(new_n708_), .C2(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n660_), .B2(new_n481_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n481_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n681_), .B2(new_n713_), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n308_), .A2(new_n311_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n359_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n566_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n615_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n255_), .A3(new_n628_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n717_), .A2(new_n508_), .A3(new_n626_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n255_), .ZN(G1332gat));
  NOR2_X1   g520(.A1(new_n717_), .A2(new_n626_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n253_), .B1(new_n722_), .B2(new_n635_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n718_), .A2(new_n253_), .A3(new_n635_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n722_), .B2(new_n645_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n718_), .A2(new_n728_), .A3(new_n645_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1334gat));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n734_), .A3(new_n481_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n722_), .A2(new_n481_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G78gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT50), .B(new_n734_), .C1(new_n722_), .C2(new_n481_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT114), .ZN(G1335gat));
  INV_X1    g540(.A(new_n717_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n690_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(G85gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n628_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n678_), .A2(new_n613_), .A3(new_n716_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n628_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n745_), .ZN(G1336gat));
  INV_X1    g548(.A(G92gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(new_n750_), .A3(new_n635_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n747_), .A2(new_n635_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n750_), .ZN(G1337gat));
  NAND4_X1  g552(.A1(new_n678_), .A2(new_n716_), .A3(new_n645_), .A4(new_n613_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G99gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G99gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n645_), .A2(new_n205_), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n756_), .A2(new_n757_), .B1(new_n743_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT116), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n761_), .ZN(new_n763_));
  OAI221_X1 g562(.A(new_n763_), .B1(new_n743_), .B2(new_n758_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  NAND4_X1  g564(.A1(new_n678_), .A2(new_n716_), .A3(new_n481_), .A4(new_n613_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n481_), .A2(new_n209_), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n768_), .A2(new_n769_), .B1(new_n743_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  OAI221_X1 g572(.A(new_n773_), .B1(new_n743_), .B2(new_n770_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NOR3_X1   g574(.A1(new_n595_), .A2(new_n613_), .A3(new_n359_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n715_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(new_n715_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n337_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n346_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(KEYINPUT117), .A3(new_n356_), .A4(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n358_), .A2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n782_), .A2(new_n356_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT117), .B1(new_n785_), .B2(new_n781_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n301_), .ZN(new_n788_));
  AND4_X1   g587(.A1(new_n203_), .A2(new_n280_), .A3(new_n287_), .A4(new_n293_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n280_), .A2(new_n287_), .A3(new_n293_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n204_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(KEYINPUT55), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n790_), .A2(new_n793_), .A3(new_n204_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n304_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT56), .B(new_n304_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n788_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n595_), .B1(new_n799_), .B2(KEYINPUT58), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(new_n788_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT118), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n788_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n277_), .A2(new_n289_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n284_), .A2(new_n286_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(KEYINPUT72), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n203_), .B1(new_n807_), .B2(new_n287_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n294_), .B1(new_n808_), .B2(new_n793_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n794_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n304_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n798_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n804_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n801_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n804_), .B(KEYINPUT58), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n595_), .A4(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n359_), .A2(new_n301_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n309_), .A2(new_n310_), .A3(new_n787_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n587_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT57), .B(new_n587_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n803_), .A2(new_n818_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n780_), .B1(new_n826_), .B2(new_n613_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n635_), .A2(new_n508_), .A3(new_n483_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n359_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(new_n613_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n780_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n828_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n824_), .A2(new_n825_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n800_), .A2(new_n802_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n613_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n833_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n828_), .B1(new_n841_), .B2(KEYINPUT59), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n840_), .B(new_n842_), .C1(new_n841_), .C2(new_n828_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n836_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n359_), .A2(G113gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT120), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n831_), .B1(new_n844_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n843_), .B(new_n312_), .C1(new_n848_), .C2(new_n830_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n715_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n830_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n830_), .B2(new_n659_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n659_), .A2(G127gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT121), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n844_), .B2(new_n857_), .ZN(G1342gat));
  INV_X1    g657(.A(new_n595_), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n836_), .A2(new_n843_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n860_), .C1(new_n835_), .C2(new_n587_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n827_), .A2(new_n587_), .A3(new_n829_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT122), .B1(new_n865_), .B2(G134gat), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n862_), .A2(new_n864_), .A3(new_n866_), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n635_), .A2(new_n508_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n482_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n359_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n312_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n870_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n834_), .A2(new_n659_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT123), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n871_), .A2(new_n880_), .A3(new_n659_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n876_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n871_), .B2(new_n659_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n827_), .A2(KEYINPUT123), .A3(new_n613_), .A4(new_n870_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n876_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1346gat));
  AOI21_X1  g686(.A(G162gat), .B1(new_n871_), .B2(new_n624_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n670_), .A2(G162gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n871_), .B2(new_n889_), .ZN(G1347gat));
  INV_X1    g689(.A(new_n840_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n628_), .A2(new_n549_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n359_), .A3(new_n645_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n551_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G169gat), .B1(new_n891_), .B2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(G169gat), .B(new_n898_), .C1(new_n891_), .C2(new_n896_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n628_), .A2(new_n483_), .A3(new_n549_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n840_), .A2(new_n903_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n904_), .A2(new_n360_), .A3(new_n510_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(G1348gat));
  INV_X1    g705(.A(new_n904_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G176gat), .B1(new_n907_), .B2(new_n312_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n827_), .A2(new_n481_), .ZN(new_n909_));
  AND4_X1   g708(.A1(G176gat), .A2(new_n892_), .A3(new_n312_), .A4(new_n645_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1349gat));
  NOR3_X1   g710(.A1(new_n904_), .A2(new_n373_), .A3(new_n613_), .ZN(new_n912_));
  INV_X1    g711(.A(G183gat), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n909_), .A2(new_n645_), .A3(new_n659_), .A4(new_n892_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n904_), .B2(new_n859_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n624_), .A2(new_n374_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n904_), .B2(new_n917_), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n892_), .A2(new_n869_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n827_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n359_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n312_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n447_), .A2(KEYINPUT126), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1353gat));
  INV_X1    g724(.A(new_n919_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n834_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  AND2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n927_), .A2(new_n613_), .A3(new_n928_), .A4(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n920_), .A2(new_n659_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n928_), .ZN(G1354gat));
  OAI21_X1  g731(.A(G218gat), .B1(new_n927_), .B2(new_n859_), .ZN(new_n933_));
  NOR4_X1   g732(.A1(new_n827_), .A2(G218gat), .A3(new_n587_), .A4(new_n919_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n920_), .B2(new_n595_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT127), .B1(new_n939_), .B2(new_n934_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n937_), .A2(new_n940_), .ZN(G1355gat));
endmodule


