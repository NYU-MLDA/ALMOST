//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  XOR2_X1   g000(.A(G120gat), .B(G148gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G176gat), .B(G204gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G230gat), .A2(G233gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT64), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT9), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(KEYINPUT9), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT10), .B(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n224_));
  INV_X1    g023(.A(new_n222_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n215_), .A2(new_n219_), .A3(new_n223_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT7), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n214_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n234_), .A3(new_n214_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n228_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G57gat), .B(G64gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n237_), .A2(KEYINPUT11), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n236_), .A2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n231_), .A2(new_n234_), .A3(new_n214_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n234_), .B1(new_n231_), .B2(new_n214_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n244_), .B(new_n227_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n210_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT66), .B(new_n210_), .C1(new_n245_), .C2(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n227_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n243_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT12), .A3(new_n248_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n258_), .A3(new_n243_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n210_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n207_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n209_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(new_n253_), .A3(new_n252_), .A4(new_n206_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT68), .B(new_n207_), .C1(new_n254_), .C2(new_n260_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n266_), .A2(new_n267_), .B1(new_n268_), .B2(KEYINPUT13), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(KEYINPUT13), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n270_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G1gat), .B(G8gat), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G15gat), .B(G22gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G1gat), .A2(G8gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT14), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n276_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n275_), .A3(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G231gat), .A2(G233gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT76), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n287_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(new_n244_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n293_));
  XOR2_X1   g092(.A(G127gat), .B(G155gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n292_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(KEYINPUT17), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n292_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n302_));
  XOR2_X1   g101(.A(G43gat), .B(G50gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(G29gat), .B(G36gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G29gat), .B(G36gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(G43gat), .B(G50gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n302_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n308_), .A3(new_n302_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT15), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(KEYINPUT15), .A3(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n255_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n236_), .A2(new_n312_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G232gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n316_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(new_n321_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G190gat), .B(G218gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G134gat), .B(G162gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT36), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n328_), .B(KEYINPUT36), .Z(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n325_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT37), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n331_), .B(KEYINPUT74), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n325_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT37), .B1(new_n336_), .B2(new_n330_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n301_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n274_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n341_));
  INV_X1    g140(.A(G134gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G127gat), .ZN(new_n343_));
  INV_X1    g142(.A(G127gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G134gat), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n343_), .A2(new_n345_), .A3(KEYINPUT87), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT87), .B1(new_n343_), .B2(new_n345_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350_));
  INV_X1    g149(.A(KEYINPUT87), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n344_), .A2(G134gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n342_), .A2(G127gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n343_), .A2(new_n345_), .A3(KEYINPUT87), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n341_), .B1(new_n349_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n350_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT88), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360_));
  INV_X1    g159(.A(G141gat), .ZN(new_n361_));
  INV_X1    g160(.A(G148gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(KEYINPUT1), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT1), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(G155gat), .A3(G162gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n375_), .A3(new_n370_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G141gat), .B(G148gat), .Z(new_n377_));
  AOI22_X1  g176(.A1(new_n369_), .A2(new_n372_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n357_), .A2(new_n359_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT100), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n349_), .B2(new_n356_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT101), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT101), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n378_), .B(new_n385_), .C1(new_n349_), .C2(new_n356_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n357_), .A2(KEYINPUT100), .A3(new_n359_), .A4(new_n379_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n382_), .A2(new_n387_), .A3(KEYINPUT4), .A4(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n380_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT102), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n389_), .A2(KEYINPUT102), .A3(new_n393_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n382_), .A2(new_n387_), .A3(new_n388_), .A4(new_n390_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n396_), .A2(new_n401_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n401_), .B1(new_n406_), .B2(new_n402_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n407_), .B2(KEYINPUT104), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n389_), .A2(KEYINPUT102), .A3(new_n393_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT102), .B1(new_n389_), .B2(new_n393_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT104), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n401_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G22gat), .B(G50gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n379_), .A2(KEYINPUT29), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT28), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n417_), .A2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n416_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n379_), .A2(KEYINPUT29), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT28), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n419_), .A3(new_n415_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G228gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(KEYINPUT89), .B2(G233gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(KEYINPUT89), .B2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(G197gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n431_));
  INV_X1    g230(.A(G204gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G197gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT90), .B1(new_n430_), .B2(G204gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT21), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G211gat), .B(G218gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT91), .B1(new_n430_), .B2(G204gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n432_), .A3(G197gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(G204gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n436_), .B(new_n437_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n437_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(KEYINPUT21), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT93), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n429_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n379_), .A2(KEYINPUT29), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n451_), .B(new_n448_), .C1(new_n449_), .C2(new_n429_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n455_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n426_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT95), .ZN(new_n461_));
  INV_X1    g260(.A(new_n426_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT94), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n463_), .A3(new_n457_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n453_), .A2(KEYINPUT94), .A3(new_n454_), .A4(new_n456_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT95), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n426_), .A2(new_n467_), .A3(new_n459_), .A4(new_n457_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n461_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT22), .B(G169gat), .Z(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(G176gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G183gat), .A2(G190gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT23), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT83), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(new_n480_), .A3(KEYINPUT23), .A4(new_n477_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n474_), .A2(KEYINPUT23), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n479_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G183gat), .A2(G190gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n473_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT25), .B(G183gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT26), .B(G190gat), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n471_), .A2(KEYINPUT24), .ZN(new_n490_));
  INV_X1    g289(.A(G169gat), .ZN(new_n491_));
  INV_X1    g290(.A(G176gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n488_), .A2(new_n489_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(KEYINPUT24), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n499_));
  INV_X1    g298(.A(new_n477_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n498_), .B(new_n499_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT23), .B1(new_n476_), .B2(new_n477_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n498_), .B1(new_n474_), .B2(KEYINPUT23), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n502_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n497_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT84), .B1(new_n487_), .B2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n503_), .A2(new_n505_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n509_), .A2(new_n494_), .A3(new_n502_), .A4(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n482_), .B1(new_n478_), .B2(KEYINPUT83), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n485_), .B1(new_n512_), .B2(new_n481_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n510_), .B(new_n511_), .C1(new_n513_), .C2(new_n473_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n448_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n448_), .ZN(new_n517_));
  OAI221_X1 g316(.A(new_n471_), .B1(G176gat), .B2(new_n472_), .C1(new_n506_), .C2(new_n485_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n495_), .B1(new_n512_), .B2(new_n481_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n494_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  AOI211_X1 g320(.A(KEYINPUT97), .B(new_n495_), .C1(new_n512_), .C2(new_n481_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n517_), .B(new_n518_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT98), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n484_), .A2(new_n496_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT97), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n520_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n494_), .A3(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n529_), .A2(KEYINPUT98), .A3(new_n517_), .A4(new_n518_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n516_), .A2(new_n525_), .A3(KEYINPUT20), .A4(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G226gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G8gat), .B(G36gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G64gat), .B(G92gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n448_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n508_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(KEYINPUT20), .A3(new_n534_), .A4(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n536_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n541_), .B1(new_n536_), .B2(new_n545_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n470_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n541_), .B(KEYINPUT105), .Z(new_n549_));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n515_), .B2(new_n448_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n535_), .B1(new_n551_), .B2(new_n523_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n543_), .A2(KEYINPUT20), .A3(new_n535_), .A4(new_n544_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n545_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n535_), .B2(new_n531_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT27), .B(new_n555_), .C1(new_n557_), .C2(new_n541_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n414_), .A2(new_n469_), .A3(new_n548_), .A4(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n412_), .B1(new_n411_), .B2(new_n401_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n407_), .A2(KEYINPUT104), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n404_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n541_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n551_), .A2(new_n523_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n534_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n566_), .B2(new_n553_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n536_), .A2(new_n545_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n390_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n382_), .A2(new_n387_), .A3(new_n388_), .A4(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT103), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n400_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n570_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n389_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n571_), .B2(new_n400_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n573_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n404_), .A2(KEYINPUT33), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n406_), .A2(new_n579_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n577_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n546_), .A2(new_n547_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n562_), .A2(new_n569_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n559_), .B1(new_n583_), .B2(new_n469_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n357_), .A2(new_n359_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n515_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT85), .B(G43gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT86), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n588_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n585_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G227gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(G15gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G71gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n221_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT30), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT31), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n589_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n592_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n592_), .B2(new_n600_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n461_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n548_), .A2(new_n605_), .A3(new_n558_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT106), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n548_), .A2(new_n605_), .A3(KEYINPUT106), .A4(new_n558_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n604_), .A2(new_n562_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n584_), .A2(new_n604_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n275_), .B1(new_n285_), .B2(new_n281_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n282_), .A2(new_n276_), .A3(new_n283_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n311_), .B(new_n310_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n311_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n284_), .B(new_n286_), .C1(new_n618_), .C2(new_n309_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n617_), .A2(new_n619_), .A3(KEYINPUT77), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT77), .B1(new_n617_), .B2(new_n619_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n614_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n314_), .A2(new_n287_), .A3(new_n315_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n619_), .A3(new_n613_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G113gat), .B(G141gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT80), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT80), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n622_), .A2(new_n630_), .A3(new_n624_), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT78), .ZN(new_n633_));
  INV_X1    g432(.A(new_n621_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n617_), .A2(new_n619_), .A3(KEYINPUT77), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n613_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n624_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n622_), .A2(KEYINPUT78), .A3(new_n624_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n627_), .B(KEYINPUT79), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n612_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n340_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n562_), .A2(KEYINPUT107), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n562_), .A2(KEYINPUT107), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n645_), .A2(G1gat), .A3(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT108), .B(KEYINPUT38), .Z(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n612_), .A2(new_n332_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n301_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n642_), .A2(new_n271_), .A3(new_n272_), .A4(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n414_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n651_), .A2(new_n652_), .A3(new_n658_), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n610_), .A2(new_n611_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n569_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n581_), .A2(new_n582_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n469_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n548_), .A2(new_n469_), .A3(new_n558_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n562_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n604_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n660_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n548_), .A2(new_n558_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n332_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n655_), .A2(new_n667_), .A3(new_n668_), .A4(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G8gat), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT109), .A3(KEYINPUT39), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT109), .B1(new_n671_), .B2(KEYINPUT39), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n671_), .B2(KEYINPUT39), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n671_), .A2(new_n675_), .A3(KEYINPUT39), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n668_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n645_), .A2(G8gat), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(new_n681_), .A3(new_n683_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  AOI21_X1  g486(.A(new_n594_), .B1(new_n656_), .B2(new_n603_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT41), .ZN(new_n689_));
  INV_X1    g488(.A(new_n645_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n594_), .A3(new_n603_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n656_), .B2(new_n469_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT42), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n690_), .A2(new_n693_), .A3(new_n469_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n669_), .A2(new_n654_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n274_), .A2(new_n612_), .A3(new_n643_), .A4(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n700_), .B2(new_n562_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n648_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G29gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n273_), .A2(new_n642_), .A3(new_n301_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n334_), .A2(new_n337_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n667_), .B2(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT43), .B(new_n707_), .C1(new_n660_), .C2(new_n666_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT44), .B(new_n705_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT113), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n612_), .B2(new_n707_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n667_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n704_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(KEYINPUT44), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n703_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(KEYINPUT112), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n722_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n701_), .B1(new_n718_), .B2(new_n724_), .ZN(G1328gat));
  NOR2_X1   g524(.A1(new_n711_), .A2(KEYINPUT113), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n716_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n668_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n721_), .A2(new_n723_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G36gat), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n700_), .A2(new_n731_), .A3(new_n668_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT115), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n732_), .B(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(KEYINPUT46), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n679_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n731_), .B1(new_n738_), .B2(new_n724_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n735_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n741_), .ZN(G1329gat));
  NAND2_X1  g541(.A1(new_n700_), .A2(new_n603_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT116), .B(G43gat), .Z(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(G43gat), .B(new_n603_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n729_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT47), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(new_n745_), .C1(new_n746_), .C2(new_n729_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n700_), .B2(new_n469_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n469_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n754_), .B2(new_n724_), .ZN(G1331gat));
  NOR4_X1   g554(.A1(new_n612_), .A2(new_n273_), .A3(new_n642_), .A4(new_n339_), .ZN(new_n756_));
  INV_X1    g555(.A(G57gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n702_), .ZN(new_n758_));
  AND4_X1   g557(.A1(new_n643_), .A2(new_n653_), .A3(new_n274_), .A4(new_n654_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n562_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n760_), .B2(new_n757_), .ZN(G1332gat));
  INV_X1    g560(.A(G64gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n759_), .B2(new_n668_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT48), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n762_), .A3(new_n668_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n759_), .B2(new_n603_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n756_), .A2(new_n767_), .A3(new_n603_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1334gat));
  INV_X1    g570(.A(G78gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n759_), .B2(new_n469_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT50), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n756_), .A2(new_n772_), .A3(new_n469_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1335gat));
  NOR4_X1   g575(.A1(new_n612_), .A2(new_n273_), .A3(new_n642_), .A4(new_n699_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n211_), .A3(new_n702_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n713_), .A2(new_n714_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n273_), .A2(new_n642_), .A3(new_n654_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n562_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n782_), .B2(new_n211_), .ZN(G1336gat));
  NAND3_X1  g582(.A1(new_n777_), .A2(new_n212_), .A3(new_n668_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n781_), .A2(new_n668_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n212_), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n777_), .A2(new_n603_), .A3(new_n217_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n781_), .A2(new_n603_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n221_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n779_), .A2(new_n469_), .A3(new_n780_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT117), .A3(G106gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT117), .B1(new_n791_), .B2(G106gat), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n795_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n777_), .A2(new_n218_), .A3(new_n469_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT53), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n794_), .A2(new_n795_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n792_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1339gat));
  AOI21_X1  g604(.A(new_n648_), .B1(new_n609_), .B2(new_n608_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n613_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n619_), .A2(new_n614_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n627_), .B1(new_n623_), .B2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n629_), .A2(new_n631_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n266_), .A2(new_n267_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n642_), .A2(new_n265_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n257_), .A2(new_n210_), .A3(new_n259_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n264_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n263_), .A2(KEYINPUT55), .A3(new_n209_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n206_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n818_), .B2(KEYINPUT56), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n260_), .B1(KEYINPUT55), .B2(new_n814_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n817_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n207_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n813_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(KEYINPUT118), .A3(new_n823_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n812_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n827_), .B2(new_n332_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT120), .B1(new_n818_), .B2(KEYINPUT56), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT56), .B(new_n207_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n822_), .A2(new_n831_), .A3(new_n823_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n810_), .A2(new_n265_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n834_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n707_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n828_), .A2(KEYINPUT57), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT119), .B(new_n840_), .C1(new_n827_), .C2(new_n332_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n654_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n271_), .A2(new_n643_), .A3(new_n272_), .A4(new_n338_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT54), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n603_), .B(new_n806_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n642_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n824_), .A2(new_n853_), .A3(new_n830_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n813_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n826_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n332_), .B1(new_n856_), .B2(new_n811_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT57), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n838_), .A2(new_n835_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n841_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n301_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n604_), .B1(new_n862_), .B2(new_n844_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n850_), .A2(new_n851_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .A4(new_n806_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n643_), .B1(new_n852_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n849_), .B1(new_n867_), .B2(new_n848_), .ZN(G1340gat));
  XOR2_X1   g667(.A(KEYINPUT122), .B(G120gat), .Z(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n273_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n847_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n273_), .B1(new_n852_), .B2(new_n866_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1341gat));
  NAND2_X1  g672(.A1(new_n654_), .A2(G127gat), .ZN(new_n874_));
  AOI211_X1 g673(.A(KEYINPUT123), .B(new_n874_), .C1(new_n852_), .C2(new_n866_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n852_), .A2(new_n866_), .B1(new_n876_), .B2(new_n874_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n847_), .A2(new_n654_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n875_), .A2(new_n344_), .B1(new_n877_), .B2(new_n878_), .ZN(G1342gat));
  AOI21_X1  g678(.A(G134gat), .B1(new_n847_), .B2(new_n332_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n852_), .A2(new_n866_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT124), .B(G134gat), .Z(new_n882_));
  NOR2_X1   g681(.A1(new_n707_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n880_), .B1(new_n881_), .B2(new_n883_), .ZN(G1343gat));
  AOI21_X1  g683(.A(new_n603_), .B1(new_n862_), .B2(new_n844_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n648_), .A2(new_n664_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n643_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n361_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n273_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n362_), .ZN(G1345gat));
  INV_X1    g690(.A(new_n887_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n654_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  OR3_X1    g694(.A1(new_n887_), .A2(G162gat), .A3(new_n669_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G162gat), .B1(new_n887_), .B2(new_n707_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1347gat));
  OAI21_X1  g697(.A(new_n603_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n648_), .A2(new_n605_), .A3(new_n668_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n899_), .A2(new_n643_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n491_), .B1(new_n905_), .B2(KEYINPUT62), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n904_), .A3(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT125), .B(new_n903_), .C1(new_n901_), .C2(new_n491_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n907_), .B(new_n908_), .C1(new_n472_), .C2(new_n902_), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n899_), .A2(new_n900_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n274_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n654_), .ZN(new_n913_));
  MUX2_X1   g712(.A(new_n488_), .B(G183gat), .S(new_n913_), .Z(G1350gat));
  NAND3_X1  g713(.A1(new_n910_), .A2(new_n489_), .A3(new_n332_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n899_), .A2(new_n707_), .A3(new_n900_), .ZN(new_n916_));
  INV_X1    g715(.A(G190gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n679_), .A2(new_n562_), .A3(new_n605_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n885_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n643_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n430_), .ZN(G1352gat));
  INV_X1    g721(.A(new_n920_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n274_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n432_), .A2(KEYINPUT126), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1353gat));
  AOI21_X1  g725(.A(new_n301_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n885_), .A2(new_n919_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT127), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n885_), .A2(new_n930_), .A3(new_n919_), .A4(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1354gat));
  OR3_X1    g733(.A1(new_n920_), .A2(G218gat), .A3(new_n669_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G218gat), .B1(new_n920_), .B2(new_n707_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1355gat));
endmodule


