//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(KEYINPUT76), .B(G15gat), .ZN(new_n202_));
  INV_X1    g001(.A(G22gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  INV_X1    g004(.A(G8gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G231gat), .A2(G233gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n212_), .B(new_n213_), .Z(new_n214_));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n217_));
  INV_X1    g016(.A(G57gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(G64gat), .ZN(new_n219_));
  INV_X1    g018(.A(G64gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(G57gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G71gat), .B(G78gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n215_), .A2(new_n223_), .A3(KEYINPUT11), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n214_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G183gat), .B(G211gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT78), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G155gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT79), .Z(new_n242_));
  AND2_X1   g041(.A1(new_n238_), .A2(new_n239_), .ZN(new_n243_));
  OR3_X1    g042(.A1(new_n232_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT6), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT6), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n247_), .A2(new_n249_), .A3(KEYINPUT66), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(new_n247_), .B2(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  INV_X1    g051(.A(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n250_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G85gat), .A2(G92gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT8), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT67), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n247_), .A2(new_n249_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n247_), .A2(new_n249_), .A3(KEYINPUT66), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n265_), .B(new_n262_), .C1(new_n270_), .C2(new_n257_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT8), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n255_), .A2(KEYINPUT69), .A3(new_n256_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n255_), .B2(new_n256_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n247_), .A2(new_n249_), .A3(KEYINPUT68), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT68), .B1(new_n247_), .B2(new_n249_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n261_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n264_), .B(new_n271_), .C1(new_n272_), .C2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT10), .B(G99gat), .Z(new_n281_));
  AOI21_X1  g080(.A(new_n270_), .B1(new_n254_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT9), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT64), .B(G92gat), .ZN(new_n284_));
  INV_X1    g083(.A(G85gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n260_), .B1(new_n259_), .B2(KEYINPUT9), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n282_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT15), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT34), .ZN(new_n299_));
  INV_X1    g098(.A(new_n295_), .ZN(new_n300_));
  OAI221_X1 g099(.A(new_n297_), .B1(KEYINPUT35), .B2(new_n299_), .C1(new_n300_), .C2(new_n292_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(KEYINPUT35), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G190gat), .B(G218gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G134gat), .B(G162gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(KEYINPUT36), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(KEYINPUT36), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n303_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT37), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n303_), .A2(new_n307_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n313_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n245_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n280_), .A2(new_n230_), .A3(new_n291_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G230gat), .A2(G233gat), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n230_), .B1(new_n280_), .B2(new_n291_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI211_X1 g127(.A(new_n328_), .B(new_n230_), .C1(new_n280_), .C2(new_n291_), .ZN(new_n329_));
  OAI22_X1  g128(.A1(new_n320_), .A2(new_n321_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT74), .ZN(new_n331_));
  INV_X1    g130(.A(new_n319_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n317_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n332_), .B1(new_n333_), .B2(new_n322_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n292_), .A2(new_n231_), .A3(new_n327_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n337_), .C1(new_n321_), .C2(new_n320_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G120gat), .B(G148gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT5), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G176gat), .B(G204gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  OR2_X1    g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT13), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(KEYINPUT13), .A3(new_n345_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n316_), .A2(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n352_), .A2(KEYINPUT80), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT24), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  MUX2_X1   g155(.A(new_n355_), .B(KEYINPUT24), .S(new_n356_), .Z(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(G190gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT25), .B(G183gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n362_), .B(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n366_), .B2(new_n363_), .ZN(new_n367_));
  OR3_X1    g166(.A1(new_n361_), .A2(KEYINPUT101), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT101), .B1(new_n361_), .B2(new_n367_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G169gat), .ZN(new_n371_));
  INV_X1    g170(.A(G176gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n354_), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(KEYINPUT102), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n362_), .A2(KEYINPUT23), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n366_), .A2(KEYINPUT23), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n362_), .B(KEYINPUT84), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n363_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(KEYINPUT85), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n375_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G204gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(G197gat), .ZN(new_n387_));
  INV_X1    g186(.A(G197gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(G204gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT21), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G211gat), .B(G218gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(KEYINPUT96), .B2(new_n387_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(KEYINPUT96), .B2(new_n387_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n390_), .B(new_n391_), .C1(new_n393_), .C2(KEYINPUT21), .ZN(new_n394_));
  INV_X1    g193(.A(new_n391_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(KEYINPUT21), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n370_), .A2(new_n385_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT103), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n405_));
  INV_X1    g204(.A(G183gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT25), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(KEYINPUT25), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n358_), .B(new_n407_), .C1(new_n408_), .C2(new_n405_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n357_), .B(new_n409_), .C1(new_n379_), .C2(new_n382_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411_));
  INV_X1    g210(.A(G169gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT22), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(KEYINPUT22), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n372_), .B(new_n413_), .C1(new_n414_), .C2(new_n411_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n354_), .B(new_n415_), .C1(new_n367_), .C2(new_n384_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  AOI211_X1 g216(.A(new_n401_), .B(new_n404_), .C1(new_n417_), .C2(new_n397_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT103), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n370_), .A2(new_n385_), .A3(new_n419_), .A4(new_n398_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n400_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n404_), .B(KEYINPUT100), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n374_), .B(KEYINPUT102), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n381_), .A2(KEYINPUT85), .B1(KEYINPUT23), .B2(new_n362_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(KEYINPUT85), .B2(new_n381_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n384_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n368_), .A2(new_n369_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n397_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT20), .B1(new_n417_), .B2(new_n397_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n423_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G8gat), .B(G36gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT18), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n421_), .A2(new_n433_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n421_), .B2(new_n433_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G1gat), .B(G29gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n446_), .B1(new_n449_), .B2(KEYINPUT1), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(new_n449_), .B2(KEYINPUT1), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n447_), .B(KEYINPUT92), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT1), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(KEYINPUT93), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(KEYINPUT3), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n457_), .B(KEYINPUT2), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n453_), .A2(new_n451_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n456_), .A2(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G127gat), .B(G134gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT90), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G113gat), .B(G120gat), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n468_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(KEYINPUT91), .A3(new_n468_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n465_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n470_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n465_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT4), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n473_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n465_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n445_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT33), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n486_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n445_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n484_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n476_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n445_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT33), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n440_), .A2(new_n488_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n361_), .A2(new_n367_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n397_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n385_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n417_), .A2(new_n397_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(KEYINPUT20), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n404_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n410_), .A2(new_n416_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n401_), .B1(new_n505_), .B2(new_n398_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n430_), .A3(new_n422_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(KEYINPUT32), .A3(new_n437_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n437_), .A2(KEYINPUT32), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n421_), .A2(new_n433_), .A3(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n489_), .A2(new_n490_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n509_), .B(new_n511_), .C1(new_n512_), .C2(new_n487_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n498_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G228gat), .A2(G233gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT98), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n397_), .B1(new_n465_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT95), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n465_), .A2(new_n518_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G22gat), .B(G50gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT28), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT94), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n518_), .A3(new_n465_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G78gat), .B(G106gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n525_), .A2(new_n529_), .A3(new_n527_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n520_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n520_), .B1(new_n533_), .B2(new_n532_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n517_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(new_n533_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n519_), .B(KEYINPUT95), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n516_), .A3(new_n534_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n514_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n512_), .A2(new_n487_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT27), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n437_), .B(KEYINPUT105), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n421_), .A2(new_n433_), .A3(new_n437_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(KEYINPUT106), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT106), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n421_), .A2(new_n433_), .A3(new_n551_), .A4(new_n437_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n546_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT27), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n542_), .B(new_n545_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n544_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G227gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT88), .ZN(new_n558_));
  INV_X1    g357(.A(G71gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G99gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(new_n478_), .Z(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT89), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n417_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT31), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n556_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT107), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n553_), .A2(new_n554_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n542_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n545_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n572_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n535_), .A2(new_n536_), .A3(new_n517_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n516_), .B1(new_n540_), .B2(new_n534_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n545_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n550_), .A2(new_n552_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT27), .ZN(new_n585_));
  INV_X1    g384(.A(new_n554_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n542_), .B1(new_n498_), .B2(new_n513_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT107), .B(new_n572_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n575_), .A2(new_n580_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n212_), .B(new_n295_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n212_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n296_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n212_), .A2(new_n295_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(KEYINPUT82), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT82), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n599_), .A2(new_n602_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT81), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n599_), .A2(KEYINPUT81), .A3(new_n602_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n352_), .A2(KEYINPUT80), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n353_), .A2(new_n590_), .A3(new_n612_), .A4(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n614_), .A2(G1gat), .A3(new_n545_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT38), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n309_), .A2(new_n312_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n590_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n245_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n619_), .A2(new_n612_), .A3(new_n351_), .A4(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n545_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n616_), .A2(new_n617_), .A3(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(new_n576_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  OR3_X1    g425(.A1(new_n614_), .A2(G8gat), .A3(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1325gat));
  OAI21_X1  g429(.A(G15gat), .B1(new_n621_), .B2(new_n572_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT41), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n614_), .A2(G15gat), .A3(new_n572_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1326gat));
  OAI21_X1  g433(.A(G22gat), .B1(new_n621_), .B2(new_n543_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n542_), .A2(new_n203_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n614_), .B2(new_n637_), .ZN(G1327gat));
  NOR3_X1   g437(.A1(new_n620_), .A2(new_n350_), .A3(new_n618_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n590_), .A2(new_n612_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n578_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n618_), .B(new_n311_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n589_), .A2(new_n580_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT107), .B1(new_n556_), .B2(new_n572_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT43), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n643_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n351_), .A2(new_n612_), .A3(new_n245_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT44), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n651_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n578_), .A2(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n642_), .B1(new_n656_), .B2(new_n657_), .ZN(G1328gat));
  XNOR2_X1  g457(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n653_), .A2(new_n655_), .A3(new_n624_), .ZN(new_n660_));
  INV_X1    g459(.A(G36gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT108), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n650_), .A2(new_n652_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n654_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n650_), .A2(KEYINPUT44), .A3(new_n652_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n576_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(G36gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n624_), .A2(G36gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n641_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT109), .B1(new_n640_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n672_), .A2(new_n674_), .A3(KEYINPUT45), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n659_), .B1(new_n669_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n659_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n679_), .C1(new_n662_), .C2(new_n668_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1329gat));
  NAND3_X1  g483(.A1(new_n656_), .A2(G43gat), .A3(new_n571_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n640_), .A2(new_n572_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(G43gat), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g487(.A1(new_n653_), .A2(new_n655_), .A3(new_n543_), .ZN(new_n689_));
  INV_X1    g488(.A(G50gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n542_), .A2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT111), .Z(new_n692_));
  OAI22_X1  g491(.A1(new_n689_), .A2(new_n690_), .B1(new_n640_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g492(.A(new_n612_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n619_), .A2(new_n694_), .A3(new_n350_), .A4(new_n620_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n545_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n590_), .A2(new_n694_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n643_), .A2(new_n351_), .A3(new_n245_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n578_), .A2(new_n218_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n695_), .B2(new_n624_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  INV_X1    g502(.A(new_n699_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n220_), .A3(new_n576_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n695_), .B2(new_n572_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n559_), .A3(new_n571_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n695_), .B2(new_n543_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n543_), .A2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n699_), .B2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n620_), .A2(new_n618_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n590_), .A2(new_n694_), .A3(new_n350_), .A4(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n285_), .A3(new_n578_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n650_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n351_), .A2(new_n620_), .A3(new_n612_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n720_), .A2(new_n545_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n723_), .B2(new_n285_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n718_), .B2(new_n576_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n720_), .A2(new_n722_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n624_), .A2(new_n284_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(G1337gat));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n650_), .A2(new_n571_), .A3(new_n721_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G99gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n281_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n717_), .A2(new_n572_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(KEYINPUT114), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n730_), .B2(G99gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n729_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT113), .B1(new_n738_), .B2(KEYINPUT114), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT115), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n739_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT51), .B1(new_n744_), .B2(new_n741_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n737_), .A2(new_n729_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(new_n748_), .ZN(G1338gat));
  NAND2_X1  g548(.A1(new_n726_), .A2(new_n542_), .ZN(new_n750_));
  OR2_X1    g549(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n254_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n717_), .A2(G106gat), .A3(new_n543_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n750_), .A2(new_n752_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n757_), .B(new_n758_), .C1(new_n751_), .C2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n751_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT53), .B1(new_n761_), .B2(new_n756_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  NAND3_X1  g562(.A1(new_n316_), .A2(new_n694_), .A3(new_n351_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n612_), .A2(new_n344_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n331_), .A2(new_n769_), .A3(new_n338_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n321_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n292_), .A2(new_n231_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n325_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n771_), .A2(new_n772_), .B1(new_n774_), .B2(new_n335_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n317_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n775_), .A2(KEYINPUT55), .B1(new_n332_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n770_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT119), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n770_), .A2(new_n777_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n343_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n770_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n780_), .B1(new_n770_), .B2(new_n777_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT56), .B(new_n343_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n768_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n596_), .A2(new_n597_), .A3(new_n593_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n602_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n606_), .A2(new_n603_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n346_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n313_), .B1(new_n788_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT57), .B1(new_n793_), .B2(KEYINPUT120), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n343_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n767_), .B1(new_n797_), .B2(new_n786_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n792_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n618_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n344_), .A2(new_n791_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n344_), .A2(new_n791_), .A3(KEYINPUT121), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT122), .B1(new_n811_), .B2(new_n643_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n797_), .A2(new_n786_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT122), .B(new_n643_), .C1(new_n813_), .C2(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n794_), .B(new_n803_), .C1(new_n812_), .C2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n766_), .B1(new_n817_), .B2(new_n245_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n577_), .A2(new_n571_), .A3(new_n578_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(G113gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n612_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(KEYINPUT123), .A3(KEYINPUT59), .ZN(new_n823_));
  OR2_X1    g622(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n824_));
  NAND2_X1  g623(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n824_), .B(new_n825_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n694_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n822_), .B1(new_n827_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n351_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n820_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n351_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n829_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n820_), .B2(new_n620_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n823_), .A2(new_n826_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n620_), .A2(G127gat), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT124), .Z(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n835_), .B2(new_n837_), .ZN(G1342gat));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n820_), .A2(new_n839_), .A3(new_n313_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n643_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n842_), .B2(new_n839_), .ZN(G1343gat));
  NOR4_X1   g642(.A1(new_n576_), .A2(new_n571_), .A3(new_n543_), .A4(new_n545_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n818_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n612_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n350_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n620_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT125), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n853_), .A3(new_n620_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1346gat));
  INV_X1    g657(.A(new_n846_), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n859_), .A2(G162gat), .A3(new_n618_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G162gat), .B1(new_n859_), .B2(new_n841_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1347gat));
  NAND3_X1  g661(.A1(new_n579_), .A2(new_n576_), .A3(new_n543_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n694_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT126), .B1(new_n818_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n802_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n643_), .B1(new_n813_), .B2(KEYINPUT58), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n815_), .A3(new_n814_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n620_), .B1(new_n870_), .B2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n867_), .B(new_n864_), .C1(new_n875_), .C2(new_n766_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n876_), .A3(G169gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n866_), .A2(new_n876_), .A3(new_n879_), .A4(G169gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(KEYINPUT62), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n877_), .A2(KEYINPUT127), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n818_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n371_), .A3(new_n864_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n883_), .A3(new_n885_), .ZN(G1348gat));
  NOR2_X1   g685(.A1(new_n818_), .A2(new_n863_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n350_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n620_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n359_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n406_), .B2(new_n890_), .ZN(G1350gat));
  NAND3_X1  g691(.A1(new_n887_), .A2(new_n358_), .A3(new_n313_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n818_), .A2(new_n841_), .A3(new_n863_), .ZN(new_n894_));
  INV_X1    g693(.A(G190gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n624_), .A2(new_n571_), .A3(new_n583_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n884_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n694_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n388_), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n351_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n386_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AND2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n898_), .A2(new_n245_), .A3(new_n903_), .A4(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n898_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n620_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n907_), .B2(new_n903_), .ZN(G1354gat));
  OR3_X1    g707(.A1(new_n898_), .A2(G218gat), .A3(new_n618_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G218gat), .B1(new_n898_), .B2(new_n841_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1355gat));
endmodule


