//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT20), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(G190gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  OR3_X1    g019(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n218_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT80), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n217_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n219_), .B(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n225_), .B(new_n227_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(G197gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT21), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(KEYINPUT89), .B2(new_n233_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G197gat), .B(G204gat), .Z(new_n244_));
  OAI21_X1  g043(.A(new_n236_), .B1(new_n244_), .B2(KEYINPUT21), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n238_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n208_), .B1(new_n232_), .B2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT78), .B(G183gat), .Z(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G190gat), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n225_), .B(new_n227_), .C1(new_n249_), .C2(new_n229_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n220_), .A2(new_n221_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n220_), .A2(KEYINPUT81), .A3(new_n221_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n227_), .A2(new_n216_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n213_), .B1(new_n211_), .B2(KEYINPUT79), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(KEYINPUT79), .B2(new_n213_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n248_), .B2(KEYINPUT25), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n250_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n247_), .B1(new_n262_), .B2(new_n246_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(KEYINPUT20), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n262_), .B2(new_n246_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT95), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n237_), .B1(new_n234_), .B2(new_n233_), .ZN(new_n272_));
  OAI211_X1 g071(.A(KEYINPUT21), .B(new_n241_), .C1(new_n244_), .C2(new_n239_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n272_), .A2(new_n273_), .B1(new_n237_), .B2(new_n235_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n231_), .A4(new_n222_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT94), .B1(new_n232_), .B2(new_n246_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n270_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n271_), .B1(new_n270_), .B2(new_n278_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n207_), .B(new_n268_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT96), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n270_), .A2(new_n278_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT95), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n270_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n287_), .A2(KEYINPUT96), .A3(new_n207_), .A4(new_n268_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n268_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n206_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n283_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT78), .B(G183gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI221_X1 g095(.A(new_n257_), .B1(KEYINPUT79), .B2(new_n213_), .C1(new_n296_), .C2(new_n259_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n297_), .A2(new_n256_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n274_), .B1(new_n298_), .B2(new_n250_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n246_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n267_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n266_), .B(new_n247_), .C1(new_n262_), .C2(new_n246_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n292_), .B1(new_n303_), .B2(new_n206_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n281_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n202_), .B1(new_n293_), .B2(new_n306_), .ZN(new_n307_));
  AOI211_X1 g106(.A(KEYINPUT102), .B(new_n305_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT1), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(KEYINPUT1), .B2(new_n314_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n312_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G155gat), .B(G162gat), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(KEYINPUT84), .A3(new_n328_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n318_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n246_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n246_), .A2(KEYINPUT87), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT88), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  OAI221_X1 g139(.A(new_n246_), .B1(KEYINPUT87), .B2(new_n340_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT90), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT91), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n343_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(KEYINPUT91), .A3(new_n343_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n318_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n332_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT84), .B1(new_n327_), .B2(new_n328_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n334_), .B(new_n352_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(KEYINPUT28), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT85), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(KEYINPUT28), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n333_), .A2(new_n357_), .A3(new_n334_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G22gat), .B(G50gat), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n359_), .A2(new_n365_), .A3(new_n363_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n367_), .A2(KEYINPUT86), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT86), .B1(new_n367_), .B2(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n351_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n367_), .A2(new_n348_), .A3(new_n368_), .A4(new_n345_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(KEYINPUT92), .A3(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G71gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G99gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G15gat), .B(G43gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT82), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n382_), .B(new_n384_), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n262_), .B(KEYINPUT30), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(KEYINPUT83), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(KEYINPUT83), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n388_), .A2(new_n385_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G127gat), .B(G134gat), .Z(new_n391_));
  XOR2_X1   g190(.A(G113gat), .B(G120gat), .Z(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT31), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OR3_X1    g194(.A1(new_n389_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G1gat), .B(G29gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT100), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT99), .B(KEYINPUT4), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n393_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n393_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(new_n405_), .B2(KEYINPUT97), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n333_), .A2(new_n411_), .A3(new_n393_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n413_), .B2(KEYINPUT4), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT98), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n413_), .A2(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n404_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n403_), .C1(new_n414_), .C2(new_n417_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n398_), .A2(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n309_), .A2(new_n377_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n305_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n371_), .A2(KEYINPUT92), .A3(new_n372_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT92), .B1(new_n371_), .B2(new_n372_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n424_), .B(new_n427_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n285_), .A2(new_n286_), .B1(new_n267_), .B2(new_n263_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(KEYINPUT101), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n301_), .A2(new_n431_), .A3(new_n302_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT101), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n423_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n420_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT33), .B(new_n404_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n414_), .A2(new_n417_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n404_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n437_), .B1(new_n444_), .B2(new_n291_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n398_), .B1(new_n430_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n426_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G43gat), .B(G50gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G29gat), .B(G36gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT69), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n453_), .A2(KEYINPUT69), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n452_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n453_), .A2(KEYINPUT69), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n454_), .A3(new_n451_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(KEYINPUT73), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT73), .B1(new_n457_), .B2(new_n459_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G15gat), .B(G22gat), .ZN(new_n463_));
  INV_X1    g262(.A(G1gat), .ZN(new_n464_));
  INV_X1    g263(.A(G8gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  NOR3_X1   g268(.A1(new_n461_), .A2(new_n462_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n457_), .A2(new_n459_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n474_), .B2(new_n460_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n450_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n469_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n457_), .A2(KEYINPUT15), .A3(new_n459_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT15), .B1(new_n457_), .B2(new_n459_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n471_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n449_), .B(KEYINPUT74), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT75), .ZN(new_n486_));
  XOR2_X1   g285(.A(G113gat), .B(G141gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT76), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G169gat), .B(G197gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n484_), .A2(KEYINPUT77), .A3(new_n486_), .A4(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n476_), .A3(new_n483_), .A4(new_n490_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT77), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n484_), .A2(new_n486_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n448_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n479_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  INV_X1    g302(.A(G106gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n381_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT7), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n503_), .A2(new_n512_), .A3(new_n381_), .A4(new_n504_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT9), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n516_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT64), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n516_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT10), .B(G99gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n511_), .B1(new_n533_), .B2(G106gat), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n514_), .A2(new_n522_), .A3(new_n518_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n524_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n457_), .A2(KEYINPUT15), .A3(new_n459_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n502_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n536_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n522_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n532_), .A2(new_n534_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n472_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n539_), .A2(new_n544_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n550_), .A2(new_n551_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT36), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n555_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n555_), .B2(new_n563_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT37), .B(new_n561_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G120gat), .B(G148gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT67), .ZN(new_n577_));
  INV_X1    g376(.A(G57gat), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(G64gat), .ZN(new_n579_));
  INV_X1    g378(.A(G64gat), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(G57gat), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(G57gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(G64gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT67), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n576_), .B1(new_n586_), .B2(KEYINPUT11), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT11), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT68), .B(new_n588_), .C1(new_n582_), .C2(new_n585_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n587_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT67), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT67), .B1(new_n583_), .B2(new_n584_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT11), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT68), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n576_), .A3(KEYINPUT11), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n597_), .A2(new_n598_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n543_), .B1(new_n593_), .B2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n592_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n590_), .A4(new_n591_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n537_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(KEYINPUT12), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n593_), .A2(new_n599_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n537_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n575_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n609_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n615_), .A2(new_n611_), .A3(new_n574_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT13), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT13), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n469_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(new_n605_), .Z(new_n623_));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(KEYINPUT17), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n628_), .B(KEYINPUT17), .Z(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n623_), .B2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n570_), .A2(new_n620_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n501_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n464_), .A3(new_n423_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n620_), .A2(new_n500_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n632_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n566_), .B1(new_n426_), .B2(new_n447_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT103), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(new_n566_), .C1(new_n426_), .C2(new_n447_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n640_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n424_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n637_), .A2(new_n647_), .ZN(G1324gat));
  NAND3_X1  g447(.A1(new_n635_), .A2(new_n465_), .A3(new_n309_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(new_n309_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n651_), .B(new_n640_), .C1(new_n642_), .C2(new_n644_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n465_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n645_), .B2(new_n309_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n650_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n642_), .A2(new_n644_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n640_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n658_), .A2(new_n653_), .A3(new_n309_), .A4(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G8gat), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(KEYINPUT39), .A3(new_n655_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n649_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT40), .B(new_n649_), .C1(new_n657_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n645_), .B2(new_n398_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT105), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n670_), .A2(KEYINPUT41), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(KEYINPUT41), .ZN(new_n672_));
  INV_X1    g471(.A(new_n398_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n634_), .A2(G15gat), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT106), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n672_), .A3(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n645_), .A2(new_n377_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(G22gat), .ZN(new_n679_));
  INV_X1    g478(.A(G22gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT42), .B(new_n680_), .C1(new_n645_), .C2(new_n377_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n377_), .A2(new_n680_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT107), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n679_), .A2(new_n681_), .B1(new_n634_), .B2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n566_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n632_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n620_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n501_), .A2(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(G29gat), .A3(new_n424_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(new_n570_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n448_), .B2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT43), .B(new_n570_), .C1(new_n426_), .C2(new_n447_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n692_), .A2(new_n638_), .A3(new_n632_), .A4(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n423_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n689_), .B1(new_n698_), .B2(G29gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT108), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n696_), .A2(new_n309_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n651_), .A2(G36gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n688_), .A2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT45), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n705_), .A3(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n696_), .A2(G43gat), .A3(new_n697_), .A4(new_n398_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n688_), .A2(new_n673_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(G43gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g513(.A1(new_n696_), .A2(G50gat), .A3(new_n697_), .A4(new_n377_), .ZN(new_n715_));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  INV_X1    g515(.A(new_n377_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n688_), .B2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1331gat));
  NOR2_X1   g518(.A1(new_n448_), .A2(new_n499_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(new_n620_), .A3(new_n639_), .A4(new_n691_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n578_), .A3(new_n423_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n499_), .A2(new_n632_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n620_), .A2(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n658_), .A2(new_n423_), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(new_n578_), .ZN(G1332gat));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n580_), .A3(new_n309_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n658_), .A2(new_n309_), .A3(new_n726_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G64gat), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n730_), .A3(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n379_), .A3(new_n398_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n658_), .A2(new_n398_), .A3(new_n726_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G71gat), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n736_), .A3(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n723_), .A2(new_n741_), .A3(new_n377_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n658_), .A2(new_n377_), .A3(new_n726_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(G78gat), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n743_), .A3(G78gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n742_), .B(KEYINPUT110), .C1(new_n745_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  INV_X1    g550(.A(new_n620_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n686_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n720_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n423_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n752_), .A2(new_n499_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n692_), .A2(new_n632_), .A3(new_n693_), .A4(new_n757_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n758_), .A2(KEYINPUT111), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(KEYINPUT111), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n423_), .A2(G85gat), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT112), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n756_), .B1(new_n761_), .B2(new_n763_), .ZN(G1336gat));
  NOR3_X1   g563(.A1(new_n754_), .A2(G92gat), .A3(new_n651_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n651_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n767_));
  INV_X1    g566(.A(G92gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT113), .B(new_n766_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1337gat));
  NOR3_X1   g572(.A1(new_n754_), .A2(new_n673_), .A3(new_n533_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n673_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n381_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT51), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n775_), .C1(new_n776_), .C2(new_n381_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n755_), .A2(new_n504_), .A3(new_n377_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G106gat), .B1(new_n758_), .B2(new_n717_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  INV_X1    g587(.A(new_n725_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n789_), .B2(new_n620_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n725_), .A2(new_n618_), .A3(new_n791_), .A4(new_n619_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n788_), .B1(new_n793_), .B2(new_n691_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT54), .B(new_n570_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n610_), .A2(KEYINPUT115), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n615_), .B2(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n615_), .A2(KEYINPUT55), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n604_), .A2(new_n614_), .A3(new_n607_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n799_), .A2(new_n801_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n574_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n574_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT116), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n574_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT116), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n616_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n482_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n477_), .A2(new_n480_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n812_), .B(new_n497_), .C1(new_n813_), .C2(new_n482_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n495_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n810_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n797_), .B1(new_n807_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n808_), .A2(new_n809_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n574_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n810_), .A4(new_n816_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n570_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n499_), .A2(new_n811_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n495_), .A2(new_n814_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n617_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n566_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT57), .B(new_n566_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n824_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n632_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n796_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n309_), .A2(new_n377_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(new_n423_), .A3(new_n398_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n499_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n833_), .A2(new_n842_), .A3(new_n632_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n833_), .B2(new_n632_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n796_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n838_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n500_), .A2(KEYINPUT119), .ZN(new_n851_));
  MUX2_X1   g650(.A(KEYINPUT119), .B(new_n851_), .S(G113gat), .Z(new_n852_));
  AOI21_X1  g651(.A(new_n841_), .B1(new_n850_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n849_), .B2(new_n752_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n847_), .A2(KEYINPUT120), .A3(new_n620_), .A4(new_n848_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(G120gat), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n752_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n840_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1341gat));
  NAND4_X1  g660(.A1(new_n847_), .A2(G127gat), .A3(new_n639_), .A4(new_n848_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863_));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n863_), .B(new_n864_), .C1(new_n839_), .C2(new_n632_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n839_), .B2(new_n632_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT122), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n862_), .A2(new_n870_), .A3(new_n865_), .A4(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n849_), .B2(new_n691_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n566_), .A2(G134gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n839_), .B2(new_n874_), .ZN(G1343gat));
  NOR3_X1   g674(.A1(new_n717_), .A2(new_n424_), .A3(new_n398_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n835_), .A2(new_n651_), .A3(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n500_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n320_), .ZN(G1344gat));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n752_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n321_), .ZN(G1345gat));
  NOR2_X1   g680(.A1(new_n877_), .A2(new_n632_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n877_), .B2(new_n691_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n566_), .A2(G162gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n877_), .B2(new_n886_), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n651_), .A2(new_n425_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n377_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n845_), .A2(new_n499_), .A3(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n845_), .A2(new_n223_), .A3(new_n499_), .A4(new_n890_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(KEYINPUT62), .B1(new_n891_), .B2(G169gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT123), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(G169gat), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n893_), .A4(new_n892_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n901_), .ZN(G1348gat));
  NAND2_X1  g701(.A1(new_n845_), .A2(new_n890_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G176gat), .B1(new_n904_), .B2(new_n620_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n794_), .A2(new_n795_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n632_), .B2(new_n833_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n377_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n889_), .A2(new_n224_), .A3(new_n752_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n905_), .B1(new_n908_), .B2(new_n909_), .ZN(G1349gat));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n639_), .A3(new_n888_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n294_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913_));
  INV_X1    g712(.A(new_n209_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n639_), .A2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n903_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n912_), .A2(new_n916_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n903_), .A2(new_n913_), .A3(new_n915_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n903_), .B2(new_n691_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n685_), .A2(new_n213_), .A3(new_n212_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n903_), .B2(new_n921_), .ZN(G1351gat));
  NAND3_X1  g721(.A1(new_n377_), .A2(new_n424_), .A3(new_n673_), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT125), .Z(new_n924_));
  NOR3_X1   g723(.A1(new_n907_), .A2(new_n651_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n499_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n620_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n639_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  AND2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(new_n930_), .B2(new_n931_), .ZN(G1354gat));
  NAND2_X1  g733(.A1(new_n570_), .A2(G218gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT126), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n925_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G218gat), .B1(new_n925_), .B2(new_n685_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939_));
  OR3_X1    g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1355gat));
endmodule


