//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_;
  XNOR2_X1  g000(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G1gat), .B(G29gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT4), .ZN(new_n208_));
  AOI22_X1  g007(.A1(KEYINPUT85), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n211_), .A2(new_n213_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n214_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n219_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(KEYINPUT82), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT82), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n218_), .A2(new_n221_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n231_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n208_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT4), .B1(new_n227_), .B2(new_n232_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n207_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n206_), .B1(new_n238_), .B2(KEYINPUT94), .ZN(new_n239_));
  INV_X1    g038(.A(new_n207_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n240_), .A3(new_n235_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT94), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n207_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G8gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G92gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT18), .B(G64gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT19), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT87), .B1(new_n251_), .B2(new_n252_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n251_), .A2(KEYINPUT87), .A3(new_n252_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n256_), .A2(KEYINPUT89), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n256_), .A2(KEYINPUT89), .ZN(new_n261_));
  OR4_X1    g060(.A1(new_n252_), .A2(new_n260_), .A3(new_n261_), .A4(new_n251_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT23), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT22), .B(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G169gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n266_), .B(new_n269_), .C1(new_n270_), .C2(new_n268_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT79), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(KEYINPUT24), .C1(new_n270_), .C2(new_n268_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n265_), .B1(new_n273_), .B2(KEYINPUT24), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n271_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n263_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(KEYINPUT80), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(new_n265_), .C1(new_n273_), .C2(KEYINPUT24), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n283_), .A2(new_n277_), .A3(new_n274_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n271_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n287_), .B2(new_n263_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n250_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n263_), .A2(new_n280_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n286_), .A2(new_n259_), .A3(new_n271_), .A4(new_n262_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(KEYINPUT20), .A3(new_n291_), .A4(new_n250_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n248_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n248_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n281_), .A2(new_n288_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n292_), .B(new_n295_), .C1(new_n296_), .C2(new_n250_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n244_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n240_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n233_), .A2(new_n207_), .A3(new_n235_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n206_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT92), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n299_), .A2(KEYINPUT92), .A3(new_n300_), .A4(new_n206_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT93), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n301_), .A2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT93), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n303_), .A2(new_n309_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n298_), .A2(new_n307_), .A3(new_n308_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n299_), .A2(new_n300_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n206_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT95), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n316_), .A3(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n301_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n248_), .A2(KEYINPUT32), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n319_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n250_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n296_), .A2(new_n321_), .ZN(new_n322_));
  AND4_X1   g121(.A1(KEYINPUT20), .A2(new_n290_), .A3(new_n321_), .A4(new_n291_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n318_), .B(new_n320_), .C1(new_n324_), .C2(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n311_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n232_), .B(KEYINPUT31), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT83), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n327_), .A2(KEYINPUT83), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  INV_X1    g129(.A(G43gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n286_), .A2(new_n271_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n286_), .B2(new_n271_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n335_), .A3(new_n332_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341_));
  INV_X1    g140(.A(G15gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n328_), .B(new_n329_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT83), .A3(new_n327_), .A4(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT28), .B(G22gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n234_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G50gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(G50gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n361_), .A3(KEYINPUT90), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n263_), .B1(new_n354_), .B2(new_n234_), .ZN(new_n368_));
  INV_X1    g167(.A(G233gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n369_), .A2(KEYINPUT86), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(KEYINPUT86), .ZN(new_n371_));
  OAI21_X1  g170(.A(G228gat), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n368_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n364_), .A2(new_n375_), .A3(new_n366_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n326_), .A2(new_n351_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n329_), .A2(new_n328_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n349_), .B2(new_n345_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n346_), .A2(new_n347_), .A3(new_n328_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n374_), .B(new_n376_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n364_), .A2(new_n375_), .A3(new_n366_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n375_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n348_), .B(new_n350_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n318_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n295_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n388_), .A2(KEYINPUT27), .A3(new_n294_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT27), .B1(new_n297_), .B2(new_n294_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n378_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G15gat), .B(G22gat), .ZN(new_n394_));
  INV_X1    g193(.A(G1gat), .ZN(new_n395_));
  INV_X1    g194(.A(G8gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT14), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G8gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(G57gat), .ZN(new_n401_));
  INV_X1    g200(.A(G64gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G57gat), .A2(G64gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G78gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT11), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(new_n409_), .A3(new_n404_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n405_), .A2(new_n407_), .A3(KEYINPUT11), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n400_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G231gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G127gat), .B(G155gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G211gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(KEYINPUT16), .B(G183gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n416_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(KEYINPUT17), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT75), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G190gat), .B(G218gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G134gat), .B(G162gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT36), .ZN(new_n430_));
  AND2_X1   g229(.A1(G85gat), .A2(G92gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G85gat), .A2(G92gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT9), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n431_), .A2(new_n433_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT10), .B(G99gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  INV_X1    g244(.A(G99gat), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n446_), .A2(KEYINPUT10), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(KEYINPUT10), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT65), .B(new_n445_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n440_), .A2(new_n441_), .A3(new_n444_), .A4(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n431_), .A2(new_n432_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n446_), .A4(new_n445_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n437_), .A2(new_n438_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT8), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(KEYINPUT8), .B(new_n451_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n450_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT71), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT15), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G29gat), .B(G36gat), .Z(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n466_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n465_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n466_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT15), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n463_), .A2(new_n464_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n464_), .B1(new_n463_), .B2(new_n476_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n469_), .A2(new_n471_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n450_), .A2(new_n461_), .A3(new_n480_), .A4(new_n462_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n479_), .A2(KEYINPUT72), .A3(new_n481_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n463_), .A2(new_n476_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT71), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n463_), .A2(new_n464_), .A3(new_n476_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(KEYINPUT72), .A3(new_n481_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n482_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n481_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G232gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT34), .ZN(new_n492_));
  NOR4_X1   g291(.A1(new_n477_), .A2(new_n478_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n484_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n430_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n477_), .A2(new_n478_), .A3(new_n490_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n483_), .B1(new_n498_), .B2(KEYINPUT72), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n488_), .A2(new_n482_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n492_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n429_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n484_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n506_), .A3(KEYINPUT74), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT73), .A3(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n507_), .A2(KEYINPUT73), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n497_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT37), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n509_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n393_), .A2(new_n426_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT64), .Z(new_n518_));
  AND2_X1   g317(.A1(new_n411_), .A2(new_n412_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n463_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n450_), .A2(new_n413_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(KEYINPUT12), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n463_), .A2(new_n523_), .A3(new_n519_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n518_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  OR3_X1    g331(.A1(new_n525_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n532_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n533_), .B(new_n534_), .C1(new_n537_), .C2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n480_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n400_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n547_), .A2(new_n400_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n476_), .A2(new_n400_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n555_), .A2(KEYINPUT76), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G169gat), .B(G197gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT77), .B(G113gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(KEYINPUT76), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n551_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT78), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n546_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n516_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n573_), .A2(KEYINPUT38), .A3(new_n395_), .A4(new_n318_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT97), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(G1gat), .B1(new_n571_), .B2(new_n572_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n577_), .A2(KEYINPUT97), .A3(KEYINPUT38), .A4(new_n318_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n568_), .A2(new_n425_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT98), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n497_), .A2(new_n506_), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n497_), .B2(new_n506_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n378_), .B2(new_n392_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(KEYINPUT98), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G1gat), .B1(new_n588_), .B2(new_n387_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT100), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n577_), .A2(new_n318_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n591_), .A2(KEYINPUT101), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT101), .B1(new_n591_), .B2(new_n592_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n579_), .B(new_n590_), .C1(new_n593_), .C2(new_n594_), .ZN(G1324gat));
  OAI21_X1  g394(.A(G8gat), .B1(new_n588_), .B2(new_n391_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT39), .ZN(new_n597_));
  INV_X1    g396(.A(new_n391_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n573_), .A2(new_n396_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n588_), .B2(new_n351_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n351_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n569_), .A2(new_n342_), .A3(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT104), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT104), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n605_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .A4(new_n611_), .ZN(G1326gat));
  OAI21_X1  g411(.A(G22gat), .B1(new_n588_), .B2(new_n377_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT42), .ZN(new_n614_));
  INV_X1    g413(.A(G22gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n377_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n569_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(G1327gat));
  AND3_X1   g417(.A1(new_n393_), .A2(KEYINPUT43), .A3(new_n514_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT43), .B1(new_n393_), .B2(new_n514_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n426_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT44), .A3(new_n568_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n393_), .A2(new_n514_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n426_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n393_), .A2(KEYINPUT43), .A3(new_n514_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n625_), .A2(new_n568_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT44), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(new_n630_), .A3(new_n318_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(G29gat), .A3(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n393_), .A2(new_n626_), .A3(new_n585_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(new_n568_), .ZN(new_n637_));
  INV_X1    g436(.A(G29gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n318_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(G1328gat));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n598_), .A2(KEYINPUT107), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n598_), .A2(KEYINPUT107), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n641_), .A3(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT45), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n630_), .A3(new_n598_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n648_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT106), .B1(new_n648_), .B2(G36gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n647_), .B(KEYINPUT46), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  NAND3_X1  g454(.A1(new_n637_), .A2(new_n331_), .A3(new_n607_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n622_), .A2(new_n607_), .A3(new_n630_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n331_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g458(.A(G50gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n616_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT108), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n637_), .A2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n622_), .A2(new_n616_), .A3(new_n630_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n660_), .ZN(G1331gat));
  INV_X1    g464(.A(new_n546_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n566_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n516_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G57gat), .B1(new_n668_), .B2(new_n318_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n586_), .A3(new_n426_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT109), .Z(new_n671_));
  NOR2_X1   g470(.A1(new_n387_), .A2(new_n401_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(G1332gat));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n402_), .A3(new_n645_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n645_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G64gat), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT48), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT48), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1333gat));
  INV_X1    g478(.A(G71gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n668_), .A2(new_n680_), .A3(new_n607_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n671_), .A2(new_n607_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(G71gat), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G71gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n668_), .A2(new_n687_), .A3(new_n616_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n671_), .A2(new_n616_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G78gat), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT50), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT50), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1335gat));
  AND2_X1   g492(.A1(new_n636_), .A2(new_n667_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G85gat), .B1(new_n694_), .B2(new_n318_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .A4(new_n667_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n318_), .A2(G85gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(G1336gat));
  AOI21_X1  g498(.A(G92gat), .B1(new_n694_), .B2(new_n598_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n645_), .A2(G92gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n697_), .B2(new_n701_), .ZN(G1337gat));
  OAI21_X1  g501(.A(G99gat), .B1(new_n696_), .B2(new_n351_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n351_), .A2(new_n443_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT111), .B1(new_n694_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g506(.A(G106gat), .B1(new_n696_), .B2(new_n377_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n710_), .B(G106gat), .C1(new_n696_), .C2(new_n377_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(KEYINPUT52), .A3(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n694_), .A2(new_n445_), .A3(new_n616_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n708_), .A2(KEYINPUT112), .A3(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g516(.A(new_n425_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n494_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n430_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT99), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n497_), .A2(new_n506_), .A3(new_n582_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n533_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT55), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n522_), .A2(new_n524_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n728_), .B(new_n729_), .C1(new_n730_), .C2(new_n518_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n518_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT55), .B1(new_n525_), .B2(KEYINPUT113), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n532_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n532_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n727_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n548_), .A2(new_n549_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n552_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n561_), .A3(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n565_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n535_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT116), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(KEYINPUT114), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n725_), .A2(new_n743_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n725_), .B2(new_n743_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n735_), .A2(new_n736_), .A3(new_n752_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n565_), .A2(new_n533_), .A3(new_n740_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n734_), .A2(new_n752_), .A3(KEYINPUT56), .A4(new_n532_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n756_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n734_), .A2(new_n532_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n532_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n758_), .B(KEYINPUT58), .C1(new_n763_), .C2(new_n752_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n514_), .A2(new_n757_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n718_), .B1(new_n750_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n507_), .A2(KEYINPUT73), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT37), .A3(new_n512_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n542_), .A2(new_n566_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n768_), .A2(new_n426_), .A3(new_n509_), .A4(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT54), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n598_), .A2(new_n387_), .A3(new_n385_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(G113gat), .A3(new_n567_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n763_), .A2(new_n727_), .B1(new_n535_), .B2(new_n741_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n719_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n746_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n725_), .A2(new_n743_), .A3(new_n747_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n514_), .A2(new_n757_), .A3(new_n764_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n626_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT117), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n786_), .A3(new_n626_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(new_n771_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n773_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n774_), .A2(KEYINPUT59), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n566_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n775_), .B1(new_n792_), .B2(G113gat), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT118), .B(new_n775_), .C1(new_n792_), .C2(G113gat), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1340gat));
  AND2_X1   g596(.A1(new_n790_), .A2(new_n791_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n774_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT119), .B(G120gat), .Z(new_n800_));
  NOR2_X1   g599(.A1(new_n666_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(KEYINPUT60), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n798_), .A2(new_n546_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n800_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(KEYINPUT60), .B2(new_n802_), .ZN(G1341gat));
  AOI21_X1  g604(.A(G127gat), .B1(new_n799_), .B2(new_n426_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n425_), .A2(G127gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n798_), .B2(new_n807_), .ZN(G1342gat));
  AOI21_X1  g607(.A(G134gat), .B1(new_n799_), .B2(new_n585_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n514_), .A2(G134gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n798_), .B2(new_n810_), .ZN(G1343gat));
  INV_X1    g610(.A(new_n382_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n770_), .B(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n425_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n812_), .B(new_n644_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT120), .B1(new_n816_), .B2(new_n387_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n382_), .B1(new_n766_), .B2(new_n771_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n318_), .A4(new_n644_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n566_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n546_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n426_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT121), .ZN(new_n827_));
  XNOR2_X1  g626(.A(KEYINPUT61), .B(G155gat), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n821_), .A2(new_n829_), .A3(new_n426_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n828_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n821_), .B2(new_n426_), .ZN(new_n833_));
  AOI211_X1 g632(.A(KEYINPUT121), .B(new_n626_), .C1(new_n817_), .C2(new_n820_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n831_), .A2(new_n835_), .ZN(G1346gat));
  AOI21_X1  g635(.A(G162gat), .B1(new_n821_), .B2(new_n585_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n514_), .A2(G162gat), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT122), .Z(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n821_), .B2(new_n839_), .ZN(G1347gat));
  NOR2_X1   g639(.A1(new_n644_), .A2(new_n318_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n607_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n616_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n788_), .A2(new_n566_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G169gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT123), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n847_), .A3(G169gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(KEYINPUT62), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(KEYINPUT123), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n267_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n849_), .B(new_n851_), .C1(new_n852_), .C2(new_n844_), .ZN(G1348gat));
  AND2_X1   g652(.A1(new_n788_), .A2(new_n843_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G176gat), .B1(new_n854_), .B2(new_n546_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n772_), .A2(new_n377_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT124), .Z(new_n857_));
  INV_X1    g656(.A(new_n842_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n666_), .A2(new_n268_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n855_), .B1(new_n859_), .B2(new_n860_), .ZN(G1349gat));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n426_), .A3(new_n858_), .ZN(new_n862_));
  INV_X1    g661(.A(G183gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n718_), .A2(new_n275_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n862_), .A2(new_n863_), .B1(new_n854_), .B2(new_n864_), .ZN(G1350gat));
  NAND2_X1  g664(.A1(new_n854_), .A2(new_n514_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G190gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n854_), .A2(new_n276_), .A3(new_n585_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1351gat));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n818_), .A2(new_n841_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n566_), .ZN(new_n872_));
  INV_X1    g671(.A(G197gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n870_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n871_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n566_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(new_n872_), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n871_), .A2(new_n546_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(G204gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT126), .B(G204gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n878_), .B2(new_n881_), .ZN(G1353gat));
  AOI21_X1  g681(.A(new_n718_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n884_), .A2(KEYINPUT127), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(KEYINPUT127), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n887_), .B(new_n888_), .Z(G1354gat));
  AOI21_X1  g688(.A(G218gat), .B1(new_n871_), .B2(new_n585_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n514_), .A2(G218gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n871_), .B2(new_n891_), .ZN(G1355gat));
endmodule


