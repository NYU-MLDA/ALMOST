//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT80), .B(G1gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G8gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT14), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT81), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n212_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT82), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n208_), .A2(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n215_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n208_), .A2(new_n212_), .A3(new_n222_), .A4(new_n216_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT83), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n217_), .A2(KEYINPUT82), .B1(new_n219_), .B2(new_n215_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n221_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n215_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n208_), .A2(new_n212_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n208_), .B2(new_n212_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n225_), .A2(new_n228_), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G169gat), .B(G197gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n225_), .A2(new_n228_), .A3(new_n234_), .A4(new_n238_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT86), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n247_), .A2(new_n244_), .A3(G183gat), .A4(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n249_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT85), .B1(new_n249_), .B2(KEYINPUT23), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n246_), .B(new_n248_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT25), .B(G183gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G190gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n253_), .B(new_n256_), .C1(new_n257_), .C2(new_n254_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT24), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(G169gat), .B2(G176gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(G169gat), .B2(G176gat), .ZN(new_n261_));
  OR3_X1    g060(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n252_), .A2(new_n258_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT87), .B(G176gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT22), .B(G169gat), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n264_), .A2(new_n265_), .B1(G169gat), .B2(G176gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n245_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n266_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT30), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT88), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G43gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(G15gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n282_), .B(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n278_), .A2(new_n280_), .A3(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G127gat), .B(G134gat), .Z(new_n288_));
  XOR2_X1   g087(.A(G113gat), .B(G120gat), .Z(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT31), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT89), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n280_), .A2(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n287_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT90), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT90), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(new_n293_), .A3(new_n292_), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n287_), .A2(new_n293_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n291_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n295_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G155gat), .ZN(new_n304_));
  INV_X1    g103(.A(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT92), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT2), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G141gat), .A3(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n311_), .A2(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT93), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT93), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n309_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n307_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n315_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n310_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n303_), .A2(KEYINPUT1), .B1(new_n304_), .B2(new_n305_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n290_), .B1(new_n321_), .B2(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n309_), .A2(new_n319_), .A3(new_n316_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n319_), .B1(new_n309_), .B2(new_n316_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n303_), .B(new_n306_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n325_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n322_), .A3(new_n310_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n290_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n327_), .A2(new_n334_), .A3(KEYINPUT4), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(new_n290_), .C1(new_n321_), .C2(new_n326_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n335_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n336_), .B(new_n341_), .C1(new_n342_), .C2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n327_), .A2(new_n334_), .A3(KEYINPUT4), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(new_n345_), .A3(new_n344_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n341_), .B1(new_n350_), .B2(new_n336_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n300_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n257_), .A2(new_n253_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n261_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT100), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n261_), .A3(KEYINPUT100), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n270_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n252_), .B1(G183gat), .B2(G190gat), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n365_), .A2(new_n367_), .B1(new_n266_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT21), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  INV_X1    g176(.A(new_n375_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n373_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n372_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n382_), .A3(new_n375_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT97), .B1(new_n378_), .B2(new_n373_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT21), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT98), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n372_), .A3(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n371_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n370_), .A2(KEYINPUT96), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT98), .B1(new_n392_), .B2(new_n385_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n381_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n369_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n381_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n387_), .B1(new_n386_), .B2(new_n372_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n392_), .A2(new_n385_), .A3(KEYINPUT98), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(new_n272_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n359_), .B1(new_n395_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n369_), .B2(new_n394_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n359_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(new_n272_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n401_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n405_), .B1(new_n401_), .B2(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n357_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n405_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n395_), .A2(new_n400_), .A3(new_n359_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n408_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n401_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT27), .A3(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(G228gat), .ZN(new_n422_));
  INV_X1    g221(.A(G233gat), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT94), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(KEYINPUT94), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT95), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT99), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n399_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n430_), .A2(new_n432_), .A3(G78gat), .ZN(new_n433_));
  INV_X1    g232(.A(G78gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n388_), .A2(new_n393_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n435_), .A2(new_n396_), .B1(new_n428_), .B2(new_n427_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT29), .B1(new_n321_), .B2(new_n326_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n421_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(G78gat), .B1(new_n430_), .B2(new_n432_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n330_), .A2(new_n332_), .A3(new_n431_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT28), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT28), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n330_), .A2(new_n332_), .A3(new_n446_), .A4(new_n431_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n427_), .A2(new_n428_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n445_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G22gat), .B(G50gat), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n321_), .A2(new_n326_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n446_), .B1(new_n455_), .B2(new_n431_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n447_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n445_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n454_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n443_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n452_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n442_), .A4(new_n439_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n420_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n355_), .A2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n364_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT100), .B1(new_n360_), .B2(new_n261_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n367_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n368_), .A2(new_n266_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n406_), .B1(new_n399_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n394_), .A2(new_n273_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n408_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n414_), .B1(new_n468_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n349_), .A2(new_n335_), .A3(new_n344_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n327_), .A2(new_n334_), .A3(new_n345_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n340_), .A3(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n477_), .A2(new_n418_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT102), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n347_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n350_), .A2(KEYINPUT102), .A3(new_n336_), .A4(new_n341_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n340_), .A2(new_n484_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n350_), .A2(new_n336_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT101), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT101), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n350_), .A2(new_n490_), .A3(new_n336_), .A4(new_n487_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n481_), .A2(new_n486_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n401_), .A2(new_n410_), .A3(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n415_), .A2(new_n416_), .ZN(new_n496_));
  OAI221_X1 g295(.A(new_n495_), .B1(new_n496_), .B2(new_n494_), .C1(new_n348_), .C2(new_n351_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n493_), .A2(new_n497_), .B1(new_n464_), .B2(new_n461_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n461_), .A2(new_n413_), .A3(new_n464_), .A4(new_n419_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(new_n353_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n300_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n467_), .B1(new_n501_), .B2(KEYINPUT104), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT104), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(new_n300_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n243_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n506_));
  OR3_X1    g305(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  INV_X1    g307(.A(G99gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n421_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G85gat), .B(G92gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT8), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT8), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n518_), .A3(new_n515_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n511_), .ZN(new_n522_));
  INV_X1    g321(.A(G85gat), .ZN(new_n523_));
  INV_X1    g322(.A(G92gat), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT9), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n521_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT65), .B(G106gat), .ZN(new_n527_));
  OR2_X1    g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n528_), .A2(KEYINPUT64), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT64), .B1(new_n528_), .B2(new_n529_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n517_), .A2(new_n519_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT11), .ZN(new_n534_));
  NAND2_X1  g333(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n536_), .A2(new_n537_), .A3(G78gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n539_));
  INV_X1    g338(.A(G71gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n434_), .B1(new_n541_), .B2(new_n535_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n534_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(G78gat), .B1(new_n536_), .B2(new_n537_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n434_), .A3(new_n535_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT11), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n544_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n549_), .A2(new_n545_), .A3(new_n546_), .A4(KEYINPUT11), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n548_), .A2(KEYINPUT67), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT67), .B1(new_n548_), .B2(new_n550_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n533_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT68), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n533_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(KEYINPUT67), .A3(new_n550_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(new_n533_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT12), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT69), .B1(new_n548_), .B2(new_n550_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n548_), .A2(KEYINPUT69), .A3(new_n550_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n533_), .A2(new_n565_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n558_), .A2(new_n565_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n553_), .A2(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n564_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n564_), .B2(new_n573_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n506_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n564_), .A2(new_n573_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n564_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT71), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n581_), .A2(new_n586_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n593_), .B2(KEYINPUT13), .ZN(new_n594_));
  AOI211_X1 g393(.A(KEYINPUT73), .B(new_n587_), .C1(new_n581_), .C2(new_n586_), .ZN(new_n595_));
  OAI22_X1  g394(.A1(new_n590_), .A2(new_n591_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT76), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT77), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT36), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n603_));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(KEYINPUT35), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(KEYINPUT35), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT75), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n608_), .B2(KEYINPUT78), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n533_), .A2(new_n215_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n556_), .A2(new_n216_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n608_), .A2(KEYINPUT78), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n615_), .A2(new_n609_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n601_), .A2(KEYINPUT36), .ZN(new_n617_));
  AND4_X1   g416(.A1(new_n602_), .A2(new_n614_), .A3(new_n616_), .A4(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n602_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT79), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT79), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n624_), .A3(new_n616_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n602_), .A2(new_n617_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n621_), .B1(new_n629_), .B2(new_n620_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n219_), .B(new_n632_), .Z(new_n633_));
  INV_X1    g432(.A(new_n569_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n635_), .A2(new_n636_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n633_), .A2(new_n634_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n551_), .A2(new_n552_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n633_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n633_), .A2(new_n644_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n640_), .B(KEYINPUT17), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n631_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n505_), .A2(new_n596_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n352_), .A2(new_n203_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT38), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n501_), .A2(KEYINPUT104), .ZN(new_n655_));
  INV_X1    g454(.A(new_n467_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n504_), .A3(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT105), .A3(new_n629_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT105), .B1(new_n657_), .B2(new_n629_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n591_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n588_), .A2(new_n589_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n593_), .A2(KEYINPUT13), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT73), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n593_), .A2(new_n592_), .A3(KEYINPUT13), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n661_), .A2(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n666_), .A2(new_n649_), .A3(new_n243_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G1gat), .B1(new_n668_), .B2(new_n352_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n654_), .A2(new_n669_), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  INV_X1    g470(.A(new_n420_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n672_), .B(new_n667_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(G8gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n673_), .B2(G8gat), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT39), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(G8gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(KEYINPUT106), .A3(new_n677_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n420_), .A2(G8gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n651_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n671_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n676_), .A2(new_n677_), .B1(new_n651_), .B2(new_n681_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n676_), .A2(new_n677_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n685_), .B(KEYINPUT40), .C1(new_n686_), .C2(new_n675_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(new_n668_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n300_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G15gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT41), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n694_), .A3(G15gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n651_), .A2(new_n284_), .A3(new_n690_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT107), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n695_), .A3(new_n697_), .ZN(G1326gat));
  INV_X1    g497(.A(G22gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n465_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n651_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n689_), .A2(new_n700_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G22gat), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT42), .B(new_n699_), .C1(new_n689_), .C2(new_n700_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(new_n629_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n649_), .A2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n666_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n505_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n353_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n649_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n666_), .A2(new_n712_), .A3(new_n243_), .ZN(new_n713_));
  AOI211_X1 g512(.A(KEYINPUT43), .B(new_n630_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n657_), .B2(new_n631_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n713_), .C1(new_n714_), .C2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n719_), .B2(KEYINPUT108), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n721_), .B(new_n713_), .C1(new_n714_), .C2(new_n716_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n718_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n353_), .A2(G29gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n711_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT46), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT110), .Z(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(G36gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n722_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n717_), .A2(new_n672_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n730_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n726_), .A2(KEYINPUT46), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n505_), .A2(new_n709_), .A3(new_n730_), .A4(new_n672_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT45), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT45), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n729_), .B1(new_n736_), .B2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n734_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n728_), .B(new_n741_), .C1(new_n744_), .C2(new_n730_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1329gat));
  INV_X1    g545(.A(G43gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n300_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n749_), .B(new_n718_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n710_), .A2(new_n690_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n747_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT111), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT47), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n723_), .A2(new_n748_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n752_), .B(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n754_), .A2(new_n759_), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n710_), .B2(new_n700_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n700_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n723_), .B2(new_n762_), .ZN(G1331gat));
  NOR3_X1   g562(.A1(new_n596_), .A2(new_n649_), .A3(new_n242_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n660_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(G57gat), .A3(new_n353_), .ZN(new_n766_));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n242_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n596_), .A2(new_n649_), .A3(new_n631_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(KEYINPUT112), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n353_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n766_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT113), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n766_), .A2(new_n778_), .A3(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1332gat));
  INV_X1    g579(.A(G64gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n771_), .A2(new_n781_), .A3(new_n672_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT48), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n765_), .A2(new_n672_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G64gat), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT48), .B(new_n781_), .C1(new_n765_), .C2(new_n672_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(G1333gat));
  NAND3_X1  g586(.A1(new_n771_), .A2(new_n540_), .A3(new_n690_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n765_), .A2(new_n690_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(G71gat), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G71gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1334gat));
  NAND3_X1  g592(.A1(new_n771_), .A2(new_n434_), .A3(new_n700_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n765_), .A2(new_n700_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(G78gat), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT50), .B(new_n434_), .C1(new_n765_), .C2(new_n700_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(G1335gat));
  NAND4_X1  g598(.A1(new_n768_), .A2(new_n707_), .A3(new_n649_), .A4(new_n666_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n523_), .A3(new_n353_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n657_), .A2(new_n631_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT43), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n657_), .A2(new_n715_), .A3(new_n631_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n712_), .A2(new_n242_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n666_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT115), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n666_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n806_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n353_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n802_), .B1(new_n815_), .B2(new_n523_), .ZN(G1336gat));
  NAND3_X1  g615(.A1(new_n801_), .A2(new_n524_), .A3(new_n672_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n672_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n819_), .B2(new_n524_), .ZN(G1337gat));
  OAI211_X1 g619(.A(new_n801_), .B(new_n690_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n806_), .A2(new_n690_), .A3(new_n812_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(new_n509_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g624(.A1(new_n801_), .A2(new_n700_), .A3(new_n527_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n806_), .A2(new_n700_), .A3(new_n812_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n827_), .A2(new_n828_), .A3(G106gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n827_), .B2(G106gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n826_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT53), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n826_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1339gat));
  NOR3_X1   g634(.A1(new_n466_), .A2(new_n352_), .A3(new_n300_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n596_), .A2(new_n243_), .A3(new_n650_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n596_), .A2(KEYINPUT54), .A3(new_n243_), .A4(new_n650_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n554_), .A2(new_n560_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n568_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n556_), .B(KEYINPUT12), .C1(new_n843_), .C2(new_n566_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n551_), .A2(new_n552_), .A3(new_n533_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(KEYINPUT12), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n563_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n848_), .B(KEYINPUT55), .C1(new_n571_), .C2(new_n572_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n583_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT56), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n583_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n854_), .A2(new_n242_), .A3(new_n585_), .A4(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n229_), .B1(new_n220_), .B2(new_n231_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n858_), .B2(new_n238_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n221_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n239_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n226_), .A2(new_n229_), .A3(new_n223_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n241_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n593_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n857_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n629_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n854_), .A2(new_n865_), .A3(new_n585_), .A4(new_n856_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n630_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n579_), .B1(new_n853_), .B2(KEYINPUT56), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(KEYINPUT58), .A3(new_n865_), .A4(new_n856_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n868_), .A2(new_n869_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n867_), .B(new_n629_), .C1(KEYINPUT118), .C2(KEYINPUT57), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n712_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n836_), .B1(new_n841_), .B2(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(G113gat), .A3(new_n243_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT59), .B(new_n836_), .C1(new_n841_), .C2(new_n877_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n243_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(G113gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n880_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT119), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n880_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1340gat));
  INV_X1    g689(.A(new_n878_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(KEYINPUT60), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT120), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n596_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n892_), .B2(new_n897_), .ZN(G1341gat));
  INV_X1    g697(.A(G127gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n891_), .A2(new_n899_), .A3(new_n712_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n649_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1342gat));
  INV_X1    g701(.A(G134gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n891_), .A2(new_n903_), .A3(new_n707_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n630_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1343gat));
  OR2_X1    g705(.A1(new_n841_), .A2(new_n877_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n907_), .A2(new_n300_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n499_), .A2(new_n352_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n242_), .A3(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n666_), .A3(new_n909_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n907_), .A2(new_n300_), .A3(new_n712_), .A4(new_n909_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT121), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n916_), .A2(KEYINPUT121), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n915_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n916_), .A2(KEYINPUT121), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n917_), .A3(new_n914_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1346gat));
  NAND2_X1  g722(.A1(new_n908_), .A2(new_n909_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G162gat), .B1(new_n924_), .B2(new_n630_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n707_), .A2(new_n305_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n926_), .ZN(G1347gat));
  NOR3_X1   g726(.A1(new_n355_), .A2(new_n700_), .A3(new_n420_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n242_), .B(new_n928_), .C1(new_n841_), .C2(new_n877_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n930_));
  AND3_X1   g729(.A1(new_n929_), .A2(G169gat), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(G169gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n907_), .A2(new_n928_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n242_), .A2(new_n265_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT123), .ZN(new_n935_));
  OAI22_X1  g734(.A1(new_n931_), .A2(new_n932_), .B1(new_n933_), .B2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  OAI221_X1 g737(.A(KEYINPUT124), .B1(new_n933_), .B2(new_n935_), .C1(new_n931_), .C2(new_n932_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1348gat));
  AND2_X1   g739(.A1(new_n907_), .A2(new_n928_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n941_), .A2(G176gat), .A3(new_n666_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n666_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n264_), .B2(new_n943_), .ZN(G1349gat));
  NOR2_X1   g743(.A1(new_n933_), .A2(new_n649_), .ZN(new_n945_));
  MUX2_X1   g744(.A(G183gat), .B(new_n253_), .S(new_n945_), .Z(G1350gat));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947_));
  INV_X1    g746(.A(G190gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n941_), .B2(new_n631_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n257_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n933_), .A2(new_n950_), .A3(new_n629_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n947_), .B1(new_n949_), .B2(new_n951_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n941_), .A2(new_n257_), .A3(new_n707_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G190gat), .B1(new_n933_), .B2(new_n630_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n953_), .A2(new_n954_), .A3(KEYINPUT125), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n955_), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n420_), .A2(new_n465_), .A3(new_n353_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n908_), .A2(new_n242_), .A3(new_n957_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g758(.A1(new_n908_), .A2(new_n666_), .A3(new_n957_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g760(.A(KEYINPUT63), .B(G211gat), .Z(new_n962_));
  AND4_X1   g761(.A1(new_n712_), .A2(new_n908_), .A3(new_n957_), .A4(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n908_), .A2(new_n712_), .A3(new_n957_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n964_), .B2(new_n965_), .ZN(G1354gat));
  NAND4_X1  g765(.A1(new_n907_), .A2(new_n300_), .A3(new_n631_), .A4(new_n957_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(G218gat), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n629_), .A2(G218gat), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n907_), .A2(new_n300_), .A3(new_n957_), .A4(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n971_), .A2(KEYINPUT126), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n968_), .A2(new_n973_), .A3(new_n970_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n972_), .A2(new_n974_), .ZN(G1355gat));
endmodule


