//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_;
  NAND2_X1  g000(.A1(G1gat), .A2(G8gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT14), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n202_), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT76), .ZN(new_n209_));
  XOR2_X1   g008(.A(G1gat), .B(G8gat), .Z(new_n210_));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n205_), .A2(new_n211_), .A3(new_n207_), .A4(new_n206_), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n210_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G231gat), .A2(G233gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n215_), .B(new_n216_), .Z(new_n217_));
  XOR2_X1   g016(.A(G71gat), .B(G78gat), .Z(new_n218_));
  XNOR2_X1  g017(.A(G57gat), .B(G64gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(KEYINPUT11), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G64gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G57gat), .ZN(new_n222_));
  INV_X1    g021(.A(G57gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G64gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT11), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(KEYINPUT69), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(new_n219_), .B2(KEYINPUT11), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n220_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(KEYINPUT69), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(new_n227_), .A3(KEYINPUT11), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n224_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n230_), .A2(new_n231_), .A3(new_n234_), .A4(new_n218_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT71), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n229_), .A2(new_n235_), .A3(KEYINPUT71), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n217_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242_));
  XOR2_X1   g041(.A(G127gat), .B(G155gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT16), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G183gat), .B(G211gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n241_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n240_), .B2(new_n217_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n236_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n217_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n217_), .A2(new_n249_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n246_), .B(KEYINPUT17), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT103), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT93), .ZN(new_n256_));
  AND2_X1   g055(.A1(G228gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G155gat), .B(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n261_), .A2(KEYINPUT89), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT89), .B1(new_n261_), .B2(new_n262_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR3_X1    g064(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n260_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G155gat), .ZN(new_n271_));
  INV_X1    g070(.A(G162gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G155gat), .A3(G162gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G141gat), .ZN(new_n278_));
  INV_X1    g077(.A(G148gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n261_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n258_), .B1(new_n270_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G197gat), .ZN(new_n283_));
  INV_X1    g082(.A(G204gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT21), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT91), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n286_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n288_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n289_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n257_), .B1(new_n282_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n286_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n292_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT91), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n302_), .A2(new_n296_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n289_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n257_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n270_), .B2(new_n281_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI211_X1 g108(.A(KEYINPUT90), .B(new_n306_), .C1(new_n270_), .C2(new_n281_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n298_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n256_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n261_), .A2(new_n262_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n261_), .A2(KEYINPUT89), .A3(new_n262_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n268_), .A2(new_n267_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n259_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n280_), .A2(new_n261_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n277_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n306_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G22gat), .B(G50gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT28), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n326_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n311_), .A2(new_n312_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n312_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT90), .B1(new_n325_), .B2(new_n306_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n307_), .A2(new_n308_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n305_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(new_n298_), .ZN(new_n336_));
  OAI22_X1  g135(.A1(new_n313_), .A2(new_n330_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n311_), .A2(new_n312_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n298_), .A3(new_n332_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n256_), .A4(new_n329_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G134gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G127gat), .ZN(new_n344_));
  INV_X1    g143(.A(G127gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G134gat), .ZN(new_n346_));
  INV_X1    g145(.A(G120gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G113gat), .ZN(new_n348_));
  INV_X1    g147(.A(G113gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G120gat), .ZN(new_n350_));
  AND4_X1   g149(.A1(new_n344_), .A2(new_n346_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n344_), .A2(new_n346_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT86), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n353_), .B(new_n358_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n354_), .B(new_n355_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n270_), .A2(new_n360_), .A3(new_n281_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n353_), .A2(new_n358_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n270_), .A2(new_n281_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n362_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n359_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G57gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n361_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n368_), .B1(new_n359_), .B2(KEYINPUT4), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n377_), .B(new_n370_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n353_), .A2(new_n358_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT31), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(KEYINPUT31), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT87), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT87), .B1(new_n383_), .B2(new_n384_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(G176gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT24), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT23), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(G183gat), .A3(G190gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  OR3_X1    g197(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n393_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT25), .B(G183gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT26), .B(G190gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT81), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G183gat), .ZN(new_n409_));
  INV_X1    g208(.A(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n398_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT22), .ZN(new_n415_));
  OAI21_X1  g214(.A(G169gat), .B1(new_n415_), .B2(KEYINPUT82), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n389_), .A3(KEYINPUT22), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n418_), .A3(new_n390_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(KEYINPUT83), .A3(new_n392_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n395_), .A2(new_n397_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT84), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT83), .B1(new_n419_), .B2(new_n392_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n408_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(G71gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G99gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G43gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT85), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n419_), .A2(new_n392_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(new_n420_), .A3(new_n414_), .A4(new_n422_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n430_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n408_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n431_), .A2(new_n434_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n434_), .B1(new_n431_), .B2(new_n440_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n386_), .B(new_n388_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n441_), .A2(new_n442_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n443_), .A2(new_n444_), .B1(new_n446_), .B2(new_n385_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n381_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G226gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT19), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n438_), .A2(new_n408_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n303_), .A2(new_n304_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n404_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n389_), .A2(KEYINPUT22), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n415_), .A2(G169gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n390_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n392_), .ZN(new_n457_));
  OAI22_X1  g256(.A1(new_n453_), .A2(new_n400_), .B1(new_n421_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT20), .B1(new_n452_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n450_), .B1(new_n451_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n297_), .A2(new_n438_), .A3(new_n408_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n450_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G8gat), .B(G36gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT18), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT100), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n461_), .A2(new_n463_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n450_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n425_), .A2(new_n452_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n458_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n462_), .B1(new_n477_), .B2(new_n297_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n464_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n470_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n473_), .B2(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT27), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT27), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n451_), .A2(new_n459_), .A3(new_n450_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n464_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(new_n470_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n475_), .A2(new_n479_), .A3(new_n485_), .A4(new_n470_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n471_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n484_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  AND4_X1   g292(.A1(new_n342_), .A2(new_n448_), .A3(new_n483_), .A4(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n381_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n480_), .A2(new_n473_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT100), .B1(new_n488_), .B2(new_n470_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n472_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n495_), .B(new_n493_), .C1(new_n498_), .C2(new_n484_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT101), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n470_), .A2(KEYINPUT32), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT98), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n488_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n460_), .B2(new_n465_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT99), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT99), .ZN(new_n507_));
  AOI211_X1 g306(.A(new_n507_), .B(new_n502_), .C1(new_n460_), .C2(new_n465_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n504_), .B(new_n381_), .C1(new_n506_), .C2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n380_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n510_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n369_), .A2(new_n377_), .A3(new_n370_), .A4(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT97), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT96), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n367_), .B1(new_n359_), .B2(KEYINPUT4), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(new_n378_), .B2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n362_), .A2(new_n366_), .A3(KEYINPUT96), .A4(new_n367_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n359_), .A2(new_n361_), .A3(new_n368_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n375_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n515_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  AOI211_X1 g323(.A(KEYINPUT97), .B(new_n522_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n514_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n480_), .A2(KEYINPUT94), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n491_), .A3(new_n490_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n509_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n342_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n483_), .A2(KEYINPUT101), .A3(new_n495_), .A4(new_n493_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n501_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n445_), .A2(new_n447_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n494_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(KEYINPUT66), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(new_n540_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n547_), .B(new_n548_), .C1(G99gat), .C2(G106gat), .ZN(new_n549_));
  INV_X1    g348(.A(G106gat), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n429_), .B(new_n550_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n543_), .A2(new_n546_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT68), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(G85gat), .ZN(new_n558_));
  INV_X1    g357(.A(G92gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n554_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT8), .B1(new_n557_), .B2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n553_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n545_), .A2(new_n540_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n552_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n557_), .A2(new_n562_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n560_), .B1(new_n570_), .B2(new_n554_), .ZN(new_n571_));
  AND2_X1   g370(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n572_));
  NOR2_X1   g371(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n554_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT65), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n550_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n543_), .A2(new_n546_), .A3(new_n581_), .ZN(new_n582_));
  OAI22_X1  g381(.A1(new_n564_), .A2(new_n569_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G29gat), .B(G36gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G43gat), .B(G50gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT15), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n567_), .A2(new_n568_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n591_), .A2(KEYINPUT8), .B1(new_n553_), .B2(new_n563_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n582_), .B1(new_n577_), .B2(new_n576_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n590_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n598_), .A2(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n590_), .A2(new_n595_), .A3(new_n604_), .A4(new_n600_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n539_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(KEYINPUT74), .A3(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(KEYINPUT36), .B2(new_n538_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n603_), .A2(KEYINPUT74), .A3(new_n605_), .A4(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n255_), .B1(new_n535_), .B2(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n500_), .A2(new_n499_), .B1(new_n529_), .B2(new_n342_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n533_), .B1(new_n614_), .B2(new_n531_), .ZN(new_n615_));
  OAI211_X1 g414(.A(KEYINPUT103), .B(new_n611_), .C1(new_n615_), .C2(new_n494_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n254_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT70), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n583_), .B2(new_n236_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n594_), .A2(KEYINPUT70), .A3(new_n249_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n594_), .A2(new_n249_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n229_), .A2(KEYINPUT71), .A3(new_n235_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT71), .B1(new_n229_), .B2(new_n235_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT12), .B1(new_n592_), .B2(new_n593_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT72), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n240_), .A2(new_n630_), .A3(KEYINPUT12), .A4(new_n583_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT12), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n594_), .B2(new_n249_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n618_), .B1(new_n594_), .B2(new_n249_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n629_), .A2(new_n631_), .A3(new_n633_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n624_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(G120gat), .B(G148gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n624_), .A2(new_n635_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT13), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n209_), .A2(new_n212_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n210_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n586_), .A2(KEYINPUT77), .A3(new_n587_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT77), .ZN(new_n654_));
  INV_X1    g453(.A(new_n587_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n584_), .A2(new_n585_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n652_), .A2(new_n653_), .A3(new_n657_), .A4(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n653_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n659_), .A2(new_n661_), .A3(KEYINPUT78), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT78), .B1(new_n659_), .B2(new_n661_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n649_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n215_), .A2(new_n589_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n661_), .A3(new_n648_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(G113gat), .B(G141gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(G169gat), .B(G197gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n664_), .A2(new_n666_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n647_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n617_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT104), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT104), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n381_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n535_), .A2(new_n675_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n254_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT37), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n611_), .A2(new_n685_), .ZN(new_n686_));
  AOI211_X1 g485(.A(KEYINPUT37), .B(new_n606_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n683_), .A2(new_n646_), .A3(new_n684_), .A4(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n381_), .B(KEYINPUT102), .Z(new_n690_));
  NOR3_X1   g489(.A1(new_n689_), .A2(G1gat), .A3(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT38), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT38), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n682_), .A2(new_n692_), .A3(new_n693_), .ZN(G1324gat));
  NAND2_X1  g493(.A1(new_n483_), .A2(new_n493_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n689_), .A2(G8gat), .A3(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n617_), .A2(new_n676_), .A3(new_n695_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G8gat), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT105), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT39), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(KEYINPUT105), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n697_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT40), .B(new_n697_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1325gat));
  OAI21_X1  g508(.A(G15gat), .B1(new_n680_), .B2(new_n534_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n712_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n689_), .A2(G15gat), .A3(new_n534_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(G1326gat));
  OR3_X1    g515(.A1(new_n689_), .A2(G22gat), .A3(new_n342_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n341_), .B1(new_n679_), .B2(new_n678_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G22gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G22gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1327gat));
  NOR3_X1   g521(.A1(new_n647_), .A2(new_n675_), .A3(new_n684_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n535_), .B2(new_n688_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n725_));
  INV_X1    g524(.A(new_n688_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(new_n726_), .C1(new_n615_), .C2(new_n494_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(KEYINPUT107), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n532_), .A2(new_n534_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n494_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n688_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n729_), .B1(new_n732_), .B2(new_n725_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n723_), .B1(new_n728_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n690_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT44), .B(new_n723_), .C1(new_n728_), .C2(new_n733_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G29gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n254_), .A2(new_n612_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT108), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n683_), .A2(new_n742_), .A3(new_n646_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n743_), .A2(KEYINPUT109), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(KEYINPUT109), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n681_), .A2(G29gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n740_), .B1(new_n746_), .B2(new_n747_), .ZN(G1328gat));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT111), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT111), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n695_), .A3(new_n738_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n736_), .A2(KEYINPUT110), .A3(new_n695_), .A4(new_n738_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(G36gat), .A3(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n696_), .A2(G36gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n744_), .A2(new_n745_), .A3(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT45), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n750_), .B(new_n751_), .C1(new_n756_), .C2(new_n759_), .ZN(new_n760_));
  AND4_X1   g559(.A1(KEYINPUT111), .A2(new_n756_), .A3(new_n749_), .A4(new_n759_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1329gat));
  NAND4_X1  g561(.A1(new_n736_), .A2(G43gat), .A3(new_n533_), .A4(new_n738_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n746_), .A2(new_n534_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(G43gat), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g565(.A(G50gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n736_), .A2(new_n341_), .A3(new_n738_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n769_), .B2(new_n768_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n341_), .A2(new_n767_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n746_), .B2(new_n772_), .ZN(G1331gat));
  INV_X1    g572(.A(new_n675_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n535_), .A2(new_n774_), .A3(new_n646_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n775_), .A2(new_n684_), .A3(new_n688_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n223_), .A3(new_n737_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n646_), .A2(new_n774_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n617_), .A2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n381_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n223_), .ZN(G1332gat));
  AOI21_X1  g580(.A(new_n221_), .B1(new_n779_), .B2(new_n695_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT48), .Z(new_n783_));
  NAND3_X1  g582(.A1(new_n776_), .A2(new_n221_), .A3(new_n695_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1333gat));
  AOI21_X1  g584(.A(new_n427_), .B1(new_n779_), .B2(new_n533_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT49), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n776_), .A2(new_n427_), .A3(new_n533_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1334gat));
  INV_X1    g588(.A(G78gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n779_), .B2(new_n341_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT50), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n776_), .A2(new_n790_), .A3(new_n341_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1335gat));
  NAND2_X1  g593(.A1(new_n775_), .A2(new_n742_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n558_), .A3(new_n737_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n728_), .A2(new_n733_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n778_), .A2(new_n254_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT113), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n381_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n797_), .B1(new_n802_), .B2(new_n558_), .ZN(G1336gat));
  NAND3_X1  g602(.A1(new_n796_), .A2(new_n559_), .A3(new_n695_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(new_n695_), .A3(new_n800_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(new_n559_), .ZN(G1337gat));
  NAND4_X1  g606(.A1(new_n796_), .A2(new_n579_), .A3(new_n580_), .A4(new_n533_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT115), .Z(new_n809_));
  NAND3_X1  g608(.A1(new_n798_), .A2(new_n533_), .A3(new_n800_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(G99gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n810_), .B2(G99gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n796_), .A2(new_n550_), .A3(new_n341_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n341_), .B(new_n800_), .C1(new_n728_), .C2(new_n733_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n550_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n820_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n816_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g624(.A1(new_n664_), .A2(new_n666_), .A3(new_n672_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n648_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n665_), .A2(new_n661_), .A3(new_n649_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n671_), .A3(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(new_n829_), .A3(KEYINPUT118), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT118), .B1(new_n826_), .B2(new_n829_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n644_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n671_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n659_), .A2(new_n661_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT78), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n659_), .A2(new_n661_), .A3(KEYINPUT78), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n836_), .B1(new_n841_), .B2(new_n648_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n835_), .B1(new_n673_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n826_), .A2(new_n829_), .A3(KEYINPUT118), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT119), .A3(new_n644_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n834_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n629_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n618_), .B1(new_n850_), .B2(new_n622_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT12), .B1(new_n583_), .B2(new_n236_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n240_), .A2(KEYINPUT12), .A3(new_n583_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(KEYINPUT72), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n854_), .A2(KEYINPUT55), .A3(new_n631_), .A4(new_n634_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n635_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n851_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n641_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(KEYINPUT56), .A3(new_n641_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n858_), .B2(new_n641_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT120), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n847_), .A2(new_n849_), .A3(new_n864_), .A4(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT119), .B1(new_n845_), .B2(new_n644_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n644_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n833_), .B(new_n869_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n864_), .B(new_n866_), .C1(new_n868_), .C2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n688_), .B1(new_n871_), .B2(new_n848_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n845_), .A2(new_n645_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n644_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(KEYINPUT117), .ZN(new_n876_));
  INV_X1    g675(.A(new_n874_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n863_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n877_), .B(KEYINPUT117), .C1(new_n878_), .C2(new_n865_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n611_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n867_), .A2(new_n872_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT57), .B(new_n611_), .C1(new_n876_), .C2(new_n880_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n684_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n688_), .A2(new_n646_), .A3(new_n675_), .A4(new_n684_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n885_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n881_), .A2(new_n882_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n868_), .A2(new_n870_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n864_), .A2(new_n866_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n848_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n726_), .A3(new_n867_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n894_), .A3(new_n884_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n254_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  INV_X1    g696(.A(new_n888_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n889_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n695_), .A2(new_n341_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n533_), .A3(new_n737_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G113gat), .B1(new_n905_), .B2(new_n774_), .ZN(new_n906_));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n902_), .C1(new_n896_), .C2(new_n898_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n904_), .B2(KEYINPUT59), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n675_), .A2(new_n349_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT123), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n906_), .B1(new_n908_), .B2(new_n910_), .ZN(G1340gat));
  OAI21_X1  g710(.A(new_n347_), .B1(new_n646_), .B2(KEYINPUT60), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n905_), .B(new_n912_), .C1(KEYINPUT60), .C2(new_n347_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n908_), .A2(new_n647_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n347_), .ZN(G1341gat));
  NAND3_X1  g714(.A1(new_n905_), .A2(new_n345_), .A3(new_n684_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n908_), .A2(new_n684_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n345_), .ZN(G1342gat));
  NAND3_X1  g717(.A1(new_n905_), .A2(new_n343_), .A3(new_n612_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n908_), .A2(new_n726_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n343_), .ZN(G1343gat));
  AOI21_X1  g720(.A(new_n533_), .B1(new_n889_), .B2(new_n899_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n695_), .A2(new_n342_), .A3(new_n690_), .ZN(new_n923_));
  AOI21_X1  g722(.A(KEYINPUT124), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n897_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n925_));
  AOI211_X1 g724(.A(KEYINPUT122), .B(new_n888_), .C1(new_n895_), .C2(new_n254_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n534_), .B(new_n923_), .C1(new_n925_), .C2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n774_), .B1(new_n924_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G141gat), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n278_), .B(new_n774_), .C1(new_n924_), .C2(new_n929_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1344gat));
  OAI21_X1  g732(.A(new_n647_), .B1(new_n924_), .B2(new_n929_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G148gat), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n279_), .B(new_n647_), .C1(new_n924_), .C2(new_n929_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1345gat));
  OAI21_X1  g736(.A(new_n684_), .B1(new_n924_), .B2(new_n929_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT61), .B(G155gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n939_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n684_), .B(new_n941_), .C1(new_n924_), .C2(new_n929_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1346gat));
  NOR2_X1   g742(.A1(new_n924_), .A2(new_n929_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n612_), .A2(new_n272_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n922_), .A2(KEYINPUT124), .A3(new_n923_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n927_), .A2(new_n928_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n688_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  OAI22_X1  g747(.A1(new_n944_), .A2(new_n945_), .B1(new_n948_), .B2(new_n272_), .ZN(G1347gat));
  NAND3_X1  g748(.A1(new_n695_), .A2(new_n533_), .A3(new_n690_), .ZN(new_n950_));
  AOI211_X1 g749(.A(new_n341_), .B(new_n950_), .C1(new_n896_), .C2(new_n898_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT125), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n952_), .A2(new_n774_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n774_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(G169gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n955_), .A2(KEYINPUT62), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n955_), .A2(KEYINPUT62), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n953_), .B1(new_n956_), .B2(new_n957_), .ZN(G1348gat));
  AOI21_X1  g757(.A(G176gat), .B1(new_n952_), .B2(new_n647_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n341_), .B1(new_n889_), .B2(new_n899_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n950_), .A2(new_n646_), .A3(new_n390_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n959_), .B1(new_n960_), .B2(new_n961_), .ZN(G1349gat));
  NOR2_X1   g761(.A1(new_n950_), .A2(new_n254_), .ZN(new_n963_));
  AOI21_X1  g762(.A(G183gat), .B1(new_n960_), .B2(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n254_), .A2(new_n402_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n952_), .B2(new_n965_), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n952_), .A2(new_n612_), .A3(new_n403_), .ZN(new_n967_));
  AND2_X1   g766(.A1(new_n952_), .A2(new_n726_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n968_), .B2(new_n410_), .ZN(G1351gat));
  AND2_X1   g768(.A1(new_n695_), .A2(new_n495_), .ZN(new_n970_));
  OAI211_X1 g769(.A(new_n534_), .B(new_n970_), .C1(new_n925_), .C2(new_n926_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n971_), .A2(new_n675_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(new_n283_), .ZN(G1352gat));
  INV_X1    g772(.A(new_n971_), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n974_), .B(new_n647_), .C1(KEYINPUT126), .C2(new_n284_), .ZN(new_n975_));
  XOR2_X1   g774(.A(KEYINPUT126), .B(G204gat), .Z(new_n976_));
  OAI21_X1  g775(.A(new_n976_), .B1(new_n971_), .B2(new_n646_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n977_), .ZN(G1353gat));
  NOR2_X1   g777(.A1(new_n971_), .A2(new_n254_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n979_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980_));
  XOR2_X1   g779(.A(KEYINPUT63), .B(G211gat), .Z(new_n981_));
  AOI21_X1  g780(.A(new_n980_), .B1(new_n979_), .B2(new_n981_), .ZN(G1354gat));
  NOR2_X1   g781(.A1(new_n611_), .A2(G218gat), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n974_), .A2(new_n983_), .ZN(new_n984_));
  OAI21_X1  g783(.A(G218gat), .B1(new_n971_), .B2(new_n688_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(KEYINPUT127), .ZN(new_n987_));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n984_), .A2(new_n988_), .A3(new_n985_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n987_), .A2(new_n989_), .ZN(G1355gat));
endmodule


