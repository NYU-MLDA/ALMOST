//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT88), .A2(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(KEYINPUT22), .C1(new_n219_), .C2(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(KEYINPUT22), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n220_), .B(new_n221_), .C1(new_n218_), .C2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .A4(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT85), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n211_), .A2(new_n212_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT25), .B(G183gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n217_), .A4(new_n228_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n231_), .B1(new_n236_), .B2(KEYINPUT86), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n224_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(G15gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT31), .ZN(new_n244_));
  INV_X1    g043(.A(new_n242_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n224_), .B(new_n245_), .C1(new_n238_), .C2(new_n237_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n208_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n247_), .A3(new_n207_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n202_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT91), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n255_), .B(new_n256_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(KEYINPUT91), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n250_), .A2(new_n252_), .A3(new_n202_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n261_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n253_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(KEYINPUT91), .ZN(new_n266_));
  INV_X1    g065(.A(new_n258_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(G155gat), .A3(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT94), .ZN(new_n273_));
  INV_X1    g072(.A(G155gat), .ZN(new_n274_));
  INV_X1    g073(.A(G162gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT93), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT1), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT93), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(G155gat), .B2(G162gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n270_), .B1(new_n273_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n268_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n269_), .B(KEYINPUT2), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n266_), .B(new_n267_), .C1(new_n283_), .C2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n273_), .A2(new_n282_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n268_), .A2(new_n269_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n293_), .A3(new_n259_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n293_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n260_), .A3(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT103), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G29gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G85gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G57gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  NAND4_X1  g106(.A1(new_n295_), .A2(KEYINPUT103), .A3(new_n297_), .A4(new_n300_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n289_), .A2(new_n294_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n296_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n303_), .A2(new_n307_), .A3(new_n308_), .A4(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n301_), .A2(new_n302_), .B1(new_n309_), .B2(new_n296_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n307_), .B1(new_n313_), .B2(new_n308_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n262_), .A2(new_n265_), .A3(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT97), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  XOR2_X1   g126(.A(KEYINPUT22), .B(G169gat), .Z(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(G176gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n217_), .B(KEYINPUT101), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n213_), .A3(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n225_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT100), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n233_), .B(KEYINPUT98), .ZN(new_n337_));
  INV_X1    g136(.A(new_n232_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n227_), .A2(new_n217_), .A3(new_n228_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n332_), .A2(new_n333_), .ZN(new_n340_));
  OAI22_X1  g139(.A1(new_n337_), .A2(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n331_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G197gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT95), .A3(G204gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT21), .B(new_n344_), .C1(new_n346_), .C2(KEYINPUT95), .ZN(new_n347_));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348_));
  INV_X1    g147(.A(KEYINPUT21), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n345_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n345_), .A2(new_n349_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n347_), .A2(new_n350_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n327_), .B1(new_n342_), .B2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n224_), .B(new_n352_), .C1(new_n238_), .C2(new_n237_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n326_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n239_), .A2(new_n353_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n352_), .B(new_n331_), .C1(new_n336_), .C2(new_n341_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT20), .A4(new_n325_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n322_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n331_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT100), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n335_), .B(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n339_), .A2(new_n340_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT98), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n233_), .B(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n367_), .B2(new_n232_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT20), .B(new_n355_), .C1(new_n369_), .C2(new_n352_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n326_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n321_), .A3(new_n359_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n361_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT106), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(KEYINPUT27), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT20), .ZN(new_n379_));
  INV_X1    g178(.A(new_n325_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n354_), .A2(new_n355_), .A3(new_n326_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n321_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n377_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n376_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT107), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G78gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G106gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G22gat), .B(G50gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT28), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n352_), .B1(new_n298_), .B2(KEYINPUT29), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n397_), .A2(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n394_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n397_), .A2(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n399_), .A3(new_n393_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n383_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n407_), .A2(KEYINPUT106), .A3(KEYINPUT27), .A4(new_n373_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n385_), .A2(new_n386_), .A3(new_n406_), .A4(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n376_), .A3(new_n384_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT107), .B1(new_n410_), .B2(new_n405_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n316_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT105), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n295_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n307_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n309_), .A2(new_n297_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n361_), .A2(new_n373_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n311_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n311_), .A2(KEYINPUT104), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT104), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n313_), .A2(new_n423_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n313_), .A2(new_n308_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n415_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n311_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n356_), .A2(new_n360_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(new_n429_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n421_), .A2(new_n425_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n413_), .B1(new_n433_), .B2(new_n405_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n314_), .B2(new_n312_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n422_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n313_), .A2(KEYINPUT33), .A3(new_n307_), .A4(new_n308_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(new_n373_), .A3(new_n361_), .A4(new_n417_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n435_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT105), .A3(new_n406_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n405_), .A2(new_n315_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n410_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n434_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n262_), .A2(new_n265_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n412_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G113gat), .B(G141gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT83), .ZN(new_n447_));
  XOR2_X1   g246(.A(G169gat), .B(G197gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G29gat), .B(G36gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G43gat), .B(G50gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n452_), .B(KEYINPUT15), .Z(new_n453_));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454_));
  INV_X1    g253(.A(G1gat), .ZN(new_n455_));
  INV_X1    g254(.A(G8gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT14), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G8gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n461_), .B2(new_n452_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n460_), .B(new_n452_), .Z(new_n466_));
  AOI22_X1  g265(.A1(new_n462_), .A2(new_n465_), .B1(new_n466_), .B2(new_n464_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n449_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT82), .B1(new_n449_), .B2(new_n470_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n467_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n445_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n390_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n479_), .A2(new_n482_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT64), .ZN(new_n486_));
  AND3_X1   g285(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT64), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n484_), .A4(new_n479_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G85gat), .B(G92gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n485_), .A2(new_n494_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(KEYINPUT8), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT65), .B(new_n495_), .C1(new_n485_), .C2(new_n494_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n494_), .A2(KEYINPUT9), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT10), .B(G99gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n390_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G85gat), .A3(G92gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n504_), .A2(new_n506_), .A3(new_n508_), .A4(new_n489_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n512_), .B2(KEYINPUT11), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n515_));
  XOR2_X1   g314(.A(G71gat), .B(G78gat), .Z(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n511_), .A3(KEYINPUT11), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(KEYINPUT11), .B2(new_n512_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n513_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT12), .B1(new_n510_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n496_), .B1(new_n486_), .B2(new_n491_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n484_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n493_), .B1(new_n528_), .B2(new_n489_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT65), .B1(new_n529_), .B2(new_n495_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n500_), .A2(new_n499_), .A3(KEYINPUT8), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n525_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT69), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n498_), .B(KEYINPUT69), .C1(new_n501_), .C2(new_n502_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n509_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT12), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n522_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n524_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n501_), .A2(new_n502_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n522_), .B(new_n509_), .C1(new_n540_), .C2(new_n525_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT70), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n541_), .A2(KEYINPUT67), .ZN(new_n549_));
  INV_X1    g348(.A(new_n509_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n523_), .B1(new_n532_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n503_), .A2(new_n552_), .A3(new_n522_), .A4(new_n509_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT68), .ZN(new_n555_));
  INV_X1    g354(.A(new_n542_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n548_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n548_), .B(KEYINPUT71), .C1(new_n557_), .C2(new_n558_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT72), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n561_), .A2(new_n569_), .A3(new_n562_), .A4(new_n566_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n548_), .B(new_n571_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT73), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n568_), .A2(KEYINPUT13), .A3(new_n570_), .A4(new_n574_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n522_), .B(new_n461_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n582_), .A2(KEYINPUT17), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT79), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT80), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n582_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n532_), .A2(new_n550_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(new_n452_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT69), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n540_), .B2(new_n525_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n550_), .B1(new_n602_), .B2(new_n534_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n603_), .B2(new_n453_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT74), .ZN(new_n608_));
  XOR2_X1   g407(.A(G134gat), .B(G162gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT36), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT76), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT75), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n606_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n595_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(new_n611_), .B2(new_n606_), .ZN(new_n618_));
  OAI22_X1  g417(.A1(new_n617_), .A2(KEYINPUT77), .B1(KEYINPUT37), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(KEYINPUT77), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n594_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n476_), .A2(new_n579_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n455_), .A3(new_n428_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT38), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n577_), .A2(new_n474_), .A3(new_n578_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT108), .ZN(new_n628_));
  INV_X1    g427(.A(new_n594_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n618_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n445_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n315_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n628_), .A2(new_n629_), .A3(new_n410_), .A4(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G8gat), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(KEYINPUT109), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT109), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n636_), .B2(G8gat), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n639_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n410_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n624_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n635_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n641_), .A2(new_n639_), .B1(new_n624_), .B2(new_n645_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n641_), .A2(new_n639_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT40), .B(new_n649_), .C1(new_n650_), .C2(new_n638_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(G1325gat));
  OAI21_X1  g451(.A(G15gat), .B1(new_n632_), .B2(new_n444_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT41), .Z(new_n654_));
  INV_X1    g453(.A(new_n444_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n624_), .A2(new_n241_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1326gat));
  XNOR2_X1  g456(.A(new_n405_), .B(KEYINPUT110), .ZN(new_n658_));
  OAI21_X1  g457(.A(G22gat), .B1(new_n632_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n658_), .A2(G22gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n623_), .B2(new_n661_), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n629_), .A2(new_n618_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n476_), .A2(new_n579_), .A3(new_n663_), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n664_), .A2(G29gat), .A3(new_n315_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n619_), .B1(KEYINPUT77), .B2(new_n617_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n410_), .A2(new_n441_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n439_), .A2(new_n406_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n413_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n655_), .B1(new_n671_), .B2(new_n440_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n667_), .B(new_n668_), .C1(new_n672_), .C2(new_n412_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n620_), .A2(new_n621_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n445_), .B2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n579_), .A2(KEYINPUT108), .A3(new_n474_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n627_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n594_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n666_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n673_), .A2(new_n675_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n682_), .A2(new_n628_), .A3(KEYINPUT44), .A4(new_n594_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(new_n428_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G29gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n665_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n644_), .A2(G36gat), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n476_), .A2(new_n579_), .A3(new_n663_), .A4(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n681_), .A2(new_n410_), .A3(new_n683_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n682_), .A2(new_n628_), .A3(new_n594_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n644_), .B1(new_n699_), .B2(new_n666_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n700_), .B2(new_n683_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT112), .B(KEYINPUT46), .C1(new_n701_), .C2(new_n693_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n697_), .A2(new_n702_), .ZN(G1329gat));
  NAND4_X1  g502(.A1(new_n681_), .A2(G43gat), .A3(new_n655_), .A4(new_n683_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n204_), .B1(new_n664_), .B2(new_n444_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g506(.A(new_n664_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n658_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G50gat), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n681_), .A2(G50gat), .A3(new_n405_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n683_), .ZN(G1331gat));
  NOR3_X1   g511(.A1(new_n579_), .A2(new_n445_), .A3(new_n474_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n622_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n428_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT113), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n579_), .A2(new_n474_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n717_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n428_), .A2(G57gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(G1332gat));
  INV_X1    g519(.A(G64gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n714_), .A2(new_n721_), .A3(new_n410_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n410_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G64gat), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT48), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT48), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n718_), .B2(new_n655_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n714_), .A2(new_n728_), .A3(new_n655_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1334gat));
  NAND3_X1  g531(.A1(new_n714_), .A2(new_n388_), .A3(new_n709_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n718_), .A2(new_n709_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G78gat), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT50), .B(new_n388_), .C1(new_n718_), .C2(new_n709_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT114), .Z(G1335gat));
  NOR3_X1   g538(.A1(new_n579_), .A2(new_n629_), .A3(new_n474_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n682_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n315_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n713_), .A2(new_n663_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n315_), .A2(G85gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n742_), .B2(new_n644_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n644_), .A2(G92gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(G1337gat));
  NAND3_X1  g549(.A1(new_n744_), .A2(new_n505_), .A3(new_n655_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n741_), .A2(new_n655_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G99gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT115), .B(new_n478_), .C1(new_n741_), .C2(new_n655_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(new_n760_));
  OAI221_X1 g559(.A(new_n751_), .B1(new_n757_), .B2(new_n758_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1338gat));
  NAND3_X1  g561(.A1(new_n744_), .A2(new_n390_), .A3(new_n405_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n741_), .A2(new_n405_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(G106gat), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT52), .B(new_n390_), .C1(new_n741_), .C2(new_n405_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n770_), .B(new_n763_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  AOI21_X1  g571(.A(new_n449_), .B1(new_n466_), .B2(new_n463_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n463_), .B1(new_n461_), .B2(new_n452_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n462_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n774_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n777_), .A2(new_n778_), .B1(new_n449_), .B2(new_n467_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT120), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n574_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n571_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n541_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n545_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n551_), .A2(new_n537_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n538_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n603_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT55), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n539_), .A2(new_n547_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n536_), .A2(new_n538_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n549_), .A2(new_n553_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n788_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n798_), .B2(new_n556_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n549_), .A2(new_n553_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n795_), .B(new_n556_), .C1(new_n790_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n794_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT118), .B(new_n794_), .C1(new_n799_), .C2(new_n802_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n784_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n571_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n808_));
  OAI22_X1  g607(.A1(KEYINPUT121), .A2(new_n807_), .B1(new_n808_), .B2(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(KEYINPUT121), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n781_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n674_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n806_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n556_), .B1(new_n790_), .B2(new_n800_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT117), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n801_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n818_), .B2(new_n794_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n783_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n810_), .C1(KEYINPUT56), .C2(new_n808_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(KEYINPUT58), .A4(new_n781_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT58), .B(new_n781_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT122), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n814_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n820_), .B1(new_n808_), .B2(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n574_), .A2(new_n474_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n575_), .A2(new_n780_), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n829_), .B(new_n630_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n566_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n805_), .A2(new_n806_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n836_), .A2(new_n782_), .B1(new_n837_), .B2(new_n783_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n834_), .B1(new_n838_), .B2(new_n831_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n839_), .B2(new_n618_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n835_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n629_), .B1(new_n828_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n622_), .A2(new_n579_), .A3(new_n475_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n842_), .A2(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n315_), .B(new_n444_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n474_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT59), .B(new_n847_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n474_), .A2(G113gat), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT123), .Z(new_n856_));
  AOI21_X1  g655(.A(new_n850_), .B1(new_n854_), .B2(new_n856_), .ZN(G1340gat));
  XNOR2_X1  g656(.A(KEYINPUT124), .B(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n579_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n849_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n579_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n858_), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n849_), .A2(new_n863_), .A3(new_n629_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n594_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n849_), .A2(new_n867_), .A3(new_n630_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n674_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1343gat));
  OR2_X1    g669(.A1(new_n842_), .A2(new_n845_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n444_), .A2(new_n405_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n315_), .A3(new_n410_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n474_), .A3(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g674(.A(new_n579_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n871_), .A2(new_n876_), .A3(new_n873_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g677(.A1(new_n871_), .A2(new_n629_), .A3(new_n873_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1346gat));
  OAI211_X1 g680(.A(new_n667_), .B(new_n873_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G162gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n618_), .A2(G162gat), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n873_), .B(new_n884_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(KEYINPUT125), .A3(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n410_), .A2(new_n315_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n444_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n474_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT126), .Z(new_n894_));
  OAI211_X1 g693(.A(new_n658_), .B(new_n894_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n895_), .A2(new_n896_), .A3(G169gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(G169gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n892_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n709_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n871_), .A2(new_n900_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n475_), .A2(new_n328_), .ZN(new_n902_));
  OAI22_X1  g701(.A1(new_n897_), .A2(new_n898_), .B1(new_n901_), .B2(new_n902_), .ZN(G1348gat));
  NAND3_X1  g702(.A1(new_n871_), .A2(new_n876_), .A3(new_n900_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n846_), .A2(new_n405_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n579_), .A2(new_n221_), .A3(new_n899_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n221_), .B1(new_n905_), .B2(new_n906_), .ZN(G1349gat));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n629_), .A3(new_n892_), .ZN(new_n908_));
  INV_X1    g707(.A(G183gat), .ZN(new_n909_));
  INV_X1    g708(.A(new_n901_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n594_), .A2(new_n367_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n908_), .A2(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1350gat));
  OAI211_X1 g711(.A(new_n667_), .B(new_n900_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G190gat), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n618_), .A2(new_n338_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n900_), .B(new_n915_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT127), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n914_), .A2(new_n919_), .A3(new_n916_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n872_), .A2(new_n891_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n871_), .A2(new_n474_), .A3(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g723(.A1(new_n871_), .A2(new_n876_), .A3(new_n922_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n871_), .A2(new_n629_), .A3(new_n922_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  NAND4_X1  g729(.A1(new_n871_), .A2(new_n629_), .A3(new_n922_), .A4(new_n930_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1354gat));
  NAND2_X1  g731(.A1(new_n871_), .A2(new_n922_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G218gat), .B1(new_n933_), .B2(new_n674_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n618_), .A2(G218gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n933_), .B2(new_n935_), .ZN(G1355gat));
endmodule


