//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT22), .B(G169gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT81), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT81), .B1(new_n210_), .B2(KEYINPUT22), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n211_), .ZN(new_n215_));
  OAI221_X1 g014(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .C1(new_n213_), .C2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT80), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n208_), .A2(KEYINPUT80), .A3(new_n219_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n225_), .B1(new_n228_), .B2(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT24), .B1(new_n210_), .B2(new_n211_), .ZN(new_n231_));
  OAI22_X1  g030(.A1(new_n226_), .A2(new_n230_), .B1(new_n217_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n222_), .B(new_n223_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n216_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G211gat), .B(G218gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(G197gat), .B(G204gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(G197gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(G197gat), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT21), .B(new_n243_), .C1(new_n247_), .C2(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n237_), .A2(KEYINPUT21), .A3(new_n247_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT90), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT21), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n238_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(new_n237_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n249_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n236_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n210_), .A2(new_n211_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n258_), .A2(new_n218_), .A3(new_n217_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n220_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n212_), .B2(new_n211_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n209_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT20), .B1(new_n265_), .B2(new_n256_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n206_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n250_), .A2(KEYINPUT90), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n254_), .A2(new_n252_), .A3(new_n237_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n268_), .A2(new_n269_), .B1(new_n240_), .B2(new_n248_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n216_), .B(new_n270_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n260_), .A2(new_n261_), .B1(new_n209_), .B2(new_n263_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n272_), .A2(new_n270_), .A3(KEYINPUT95), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT95), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n265_), .B2(new_n256_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT20), .B(new_n271_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n267_), .B1(new_n276_), .B2(new_n206_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G8gat), .B(G36gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT18), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n273_), .A2(new_n275_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(KEYINPUT20), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n206_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n266_), .B1(new_n236_), .B2(new_n256_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n205_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n288_), .A3(new_n281_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(KEYINPUT27), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT98), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n286_), .A2(new_n288_), .A3(new_n281_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n281_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n295_), .B2(KEYINPUT27), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n286_), .A2(new_n288_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n282_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n289_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT98), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n291_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n304_), .A2(new_n305_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n304_), .A2(new_n305_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n303_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n306_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(KEYINPUT85), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n303_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n315_));
  AND2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT86), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n318_), .B1(new_n324_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n318_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n320_), .A2(new_n322_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n325_), .B1(new_n316_), .B2(KEYINPUT1), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n313_), .A2(new_n315_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(new_n336_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT4), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n313_), .A2(new_n315_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n338_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n339_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G85gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT0), .B(G57gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n347_), .A2(new_n350_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT87), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OR3_X1    g163(.A1(new_n270_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n270_), .B2(new_n361_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT91), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n365_), .A2(new_n366_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(KEYINPUT92), .A3(new_n369_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n338_), .A2(KEYINPUT29), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT28), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT93), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT93), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n376_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n382_), .A2(new_n371_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n374_), .A2(new_n367_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n359_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT96), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n356_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n357_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT33), .B1(new_n395_), .B2(KEYINPUT96), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n342_), .A2(new_n348_), .A3(new_n346_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n340_), .A2(new_n344_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n357_), .B(new_n397_), .C1(new_n398_), .C2(new_n346_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n295_), .A2(new_n394_), .A3(new_n396_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n281_), .A2(KEYINPUT32), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n297_), .B2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n286_), .A2(new_n288_), .A3(KEYINPUT97), .A4(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n356_), .A2(new_n358_), .B1(new_n277_), .B2(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n400_), .A2(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n376_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n385_), .B1(new_n376_), .B2(new_n382_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n390_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n302_), .A2(new_n391_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT83), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n236_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT31), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(G71gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G99gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(new_n341_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n419_), .B(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n202_), .B1(new_n414_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n427_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT98), .B1(new_n299_), .B2(new_n300_), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n292_), .B(KEYINPUT27), .C1(new_n298_), .C2(new_n289_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n290_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n359_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n412_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n412_), .B1(new_n400_), .B2(new_n408_), .ZN(new_n436_));
  OAI211_X1 g235(.A(KEYINPUT99), .B(new_n429_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n432_), .A2(new_n412_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n429_), .A2(new_n359_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n428_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G85gat), .ZN(new_n447_));
  INV_X1    g246(.A(G92gat), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT9), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G85gat), .B(G92gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT9), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT10), .B(G99gat), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT64), .B(G106gat), .Z(new_n455_));
  OAI211_X1 g254(.A(new_n450_), .B(new_n452_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT7), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(KEYINPUT65), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(KEYINPUT7), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n459_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(KEYINPUT7), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n458_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n457_), .B(new_n451_), .C1(new_n467_), .C2(new_n446_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT66), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n442_), .A2(G99gat), .A3(G106gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT66), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n470_), .A2(new_n473_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n457_), .B1(new_n474_), .B2(new_n451_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n468_), .B1(new_n475_), .B2(KEYINPUT67), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  AOI211_X1 g276(.A(new_n477_), .B(new_n457_), .C1(new_n474_), .C2(new_n451_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n456_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G29gat), .B(G36gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT15), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT73), .ZN(new_n485_));
  INV_X1    g284(.A(new_n479_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G232gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT34), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n486_), .A2(new_n482_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n487_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G190gat), .B(G218gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT36), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(KEYINPUT36), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n494_), .A2(new_n502_), .A3(new_n495_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT100), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n441_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT68), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G71gat), .B(G78gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n510_), .B(KEYINPUT68), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT69), .B1(new_n479_), .B2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n456_), .B(new_n520_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n479_), .A2(KEYINPUT69), .A3(new_n521_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n508_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT70), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(KEYINPUT12), .ZN(new_n529_));
  INV_X1    g328(.A(new_n451_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT66), .B1(new_n471_), .B2(new_n472_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n460_), .A2(KEYINPUT65), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n458_), .B1(new_n465_), .B2(new_n532_), .ZN(new_n533_));
  AOI211_X1 g332(.A(G99gat), .B(G106gat), .C1(new_n462_), .C2(KEYINPUT7), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n530_), .B1(new_n535_), .B2(new_n473_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n477_), .B1(new_n536_), .B2(new_n457_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n475_), .A2(KEYINPUT67), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n468_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n520_), .B1(new_n539_), .B2(new_n456_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n529_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n479_), .A2(new_n542_), .A3(new_n521_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n507_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n508_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G120gat), .B(G148gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  NAND4_X1  g351(.A1(new_n528_), .A2(new_n545_), .A3(new_n547_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT72), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n547_), .A2(new_n545_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n528_), .A4(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n528_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n552_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n558_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT13), .B1(new_n558_), .B2(new_n561_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565_));
  INV_X1    g364(.A(G1gat), .ZN(new_n566_));
  INV_X1    g365(.A(G8gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G8gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n520_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT16), .ZN(new_n577_));
  XOR2_X1   g376(.A(G183gat), .B(G211gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(KEYINPUT17), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n574_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G169gat), .B(G197gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n483_), .A2(new_n571_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT75), .ZN(new_n588_));
  INV_X1    g387(.A(new_n571_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n482_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n588_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n571_), .B(new_n482_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n591_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n586_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(new_n585_), .C1(new_n594_), .C2(new_n591_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(KEYINPUT76), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n600_), .B(new_n586_), .C1(new_n592_), .C2(new_n595_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n564_), .A2(new_n582_), .A3(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n506_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n506_), .A2(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT101), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n433_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT102), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n504_), .A2(KEYINPUT37), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n501_), .A2(new_n614_), .A3(new_n503_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n582_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT74), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n562_), .A2(new_n563_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n602_), .B(KEYINPUT77), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n619_), .A2(new_n441_), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n566_), .A3(new_n359_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT38), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n612_), .A2(new_n625_), .ZN(G1324gat));
  OAI21_X1  g425(.A(G8gat), .B1(new_n605_), .B2(new_n302_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT39), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n567_), .A3(new_n432_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(G1325gat));
  INV_X1    g431(.A(G15gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n623_), .A2(new_n633_), .A3(new_n427_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n429_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n633_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(KEYINPUT41), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n635_), .A2(new_n638_), .A3(new_n633_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT104), .B(new_n634_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1326gat));
  OAI21_X1  g443(.A(G22gat), .B1(new_n610_), .B2(new_n413_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n623_), .A2(new_n647_), .A3(new_n412_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n504_), .A2(new_n582_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n622_), .A2(new_n441_), .A3(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT107), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT107), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n359_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n564_), .A2(new_n617_), .A3(new_n603_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n441_), .A2(new_n658_), .A3(new_n616_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n441_), .B2(new_n616_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n657_), .B(KEYINPUT44), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT106), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n441_), .A2(new_n616_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n441_), .A2(new_n616_), .A3(new_n658_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(KEYINPUT44), .A4(new_n657_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n662_), .A2(new_n668_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n359_), .A2(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n655_), .B1(new_n671_), .B2(new_n672_), .ZN(G1328gat));
  NOR2_X1   g472(.A1(new_n302_), .A2(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n652_), .A2(new_n653_), .A3(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n302_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n656_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n667_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n661_), .A2(KEYINPUT106), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT108), .B(new_n677_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n662_), .A2(new_n668_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT108), .B1(new_n683_), .B2(new_n677_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n676_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n676_), .B(new_n686_), .C1(new_n682_), .C2(new_n684_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  NAND2_X1  g489(.A1(new_n654_), .A2(new_n427_), .ZN(new_n691_));
  INV_X1    g490(.A(G43gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n671_), .A2(G43gat), .A3(new_n427_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n695_), .B(new_n697_), .ZN(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n654_), .B2(new_n412_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n412_), .A2(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n671_), .B2(new_n700_), .ZN(G1331gat));
  INV_X1    g500(.A(new_n506_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n620_), .A2(new_n582_), .A3(new_n621_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n702_), .A2(G57gat), .A3(new_n359_), .A4(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n564_), .A2(new_n603_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n441_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n619_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n708_), .B2(new_n433_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n704_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT112), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n704_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1332gat));
  NAND2_X1  g516(.A1(new_n702_), .A2(new_n703_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G64gat), .B1(new_n718_), .B2(new_n302_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT48), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n302_), .A2(G64gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n708_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT113), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n718_), .B2(new_n429_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n427_), .A2(new_n421_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n708_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n718_), .B2(new_n413_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n413_), .A2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n708_), .B2(new_n730_), .ZN(G1335gat));
  AND2_X1   g530(.A1(new_n707_), .A2(new_n650_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n447_), .A3(new_n359_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n666_), .A2(new_n617_), .A3(new_n706_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n359_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n736_), .B2(new_n447_), .ZN(G1336gat));
  AOI21_X1  g536(.A(new_n448_), .B1(new_n734_), .B2(new_n432_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n302_), .A2(G92gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n732_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT114), .Z(G1337gat));
  XNOR2_X1  g540(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n666_), .A2(new_n427_), .A3(new_n617_), .A4(new_n706_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G99gat), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT115), .B1(new_n743_), .B2(G99gat), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n732_), .A2(new_n453_), .A3(new_n427_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n742_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n749_), .B(new_n742_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  NOR2_X1   g552(.A1(new_n413_), .A2(new_n455_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n732_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT117), .Z(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n666_), .A2(new_n412_), .A3(new_n617_), .A4(new_n706_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(G106gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT118), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(KEYINPUT52), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n756_), .A2(new_n762_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n762_), .A2(new_n756_), .A3(new_n766_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  NAND3_X1  g570(.A1(new_n618_), .A2(new_n564_), .A3(new_n621_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n479_), .A2(new_n521_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT12), .A3(new_n523_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n508_), .A3(new_n543_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT121), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n776_), .A2(new_n779_), .A3(new_n508_), .A4(new_n543_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n776_), .A2(new_n543_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT55), .B1(new_n782_), .B2(new_n507_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n508_), .C1(new_n776_), .C2(new_n543_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n552_), .B1(new_n781_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT56), .ZN(new_n788_));
  INV_X1    g587(.A(new_n598_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n588_), .A2(G229gat), .A3(G233gat), .A4(new_n590_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n585_), .B1(new_n593_), .B2(new_n591_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(new_n558_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n558_), .A4(new_n792_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n616_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n504_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n558_), .A2(new_n603_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n602_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT120), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n787_), .B2(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n545_), .A2(new_n784_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n782_), .A2(KEYINPUT55), .A3(new_n507_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n778_), .A4(new_n780_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n560_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT122), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n560_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n803_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n558_), .A2(new_n561_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n792_), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT57), .B(new_n798_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n809_), .B2(KEYINPUT122), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n804_), .B(KEYINPUT56), .C1(new_n808_), .C2(new_n560_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n818_), .A2(new_n819_), .B1(new_n802_), .B2(KEYINPUT120), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n802_), .A2(KEYINPUT120), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n817_), .B1(new_n822_), .B2(new_n504_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n797_), .B1(new_n816_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n617_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n774_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n429_), .A2(new_n433_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n438_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n438_), .A2(new_n828_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT123), .B(new_n797_), .C1(new_n816_), .C2(new_n823_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n617_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n830_), .B1(new_n834_), .B2(new_n774_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n829_), .B1(new_n835_), .B2(new_n827_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n621_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n835_), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n838_), .A2(G113gat), .A3(new_n602_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1340gat));
  XNOR2_X1  g639(.A(KEYINPUT124), .B(G120gat), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n836_), .B2(new_n564_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n564_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n835_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n836_), .B2(new_n617_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n838_), .A2(G127gat), .A3(new_n617_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1342gat));
  INV_X1    g648(.A(new_n616_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G134gat), .B1(new_n836_), .B2(new_n850_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n838_), .A2(G134gat), .A3(new_n505_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1343gat));
  NOR4_X1   g652(.A1(new_n432_), .A2(new_n413_), .A3(new_n433_), .A4(new_n427_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n834_), .B2(new_n774_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n603_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n620_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n856_), .B2(new_n582_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n773_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n772_), .B(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n582_), .B1(new_n824_), .B2(new_n831_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n833_), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n868_), .A2(KEYINPUT125), .A3(new_n617_), .A4(new_n855_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(new_n864_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n834_), .A2(new_n774_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n582_), .A3(new_n854_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT125), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n856_), .A2(new_n863_), .A3(new_n582_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n861_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n875_), .ZN(G1346gat));
  INV_X1    g675(.A(new_n856_), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n877_), .A2(G162gat), .A3(new_n505_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G162gat), .B1(new_n877_), .B2(new_n850_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1347gat));
  NAND2_X1  g679(.A1(new_n439_), .A2(new_n432_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n412_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n826_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883_), .B2(new_n602_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n885_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n883_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n212_), .A3(new_n603_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n887_), .A3(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(G176gat), .B1(new_n888_), .B2(new_n620_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n868_), .A2(new_n412_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n564_), .A2(new_n211_), .A3(new_n881_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n883_), .A2(new_n227_), .A3(new_n617_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n892_), .A2(new_n432_), .A3(new_n439_), .A4(new_n582_), .ZN(new_n896_));
  INV_X1    g695(.A(G183gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n883_), .B2(new_n850_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n505_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n224_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n883_), .B2(new_n901_), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n302_), .A2(new_n434_), .A3(new_n427_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n868_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n603_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n620_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g708(.A1(new_n871_), .A2(new_n903_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT63), .B(G211gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n617_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n905_), .A2(new_n582_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  NOR3_X1   g714(.A1(new_n868_), .A2(new_n505_), .A3(new_n904_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G218gat), .B1(new_n916_), .B2(KEYINPUT126), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n910_), .B2(new_n505_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n616_), .A2(G218gat), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT127), .Z(new_n921_));
  AOI22_X1  g720(.A1(new_n917_), .A2(new_n919_), .B1(new_n905_), .B2(new_n921_), .ZN(G1355gat));
endmodule


