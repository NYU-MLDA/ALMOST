//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n973_, new_n974_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_,
    new_n995_, new_n996_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT91), .B1(new_n204_), .B2(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT91), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(G197gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  INV_X1    g010(.A(G218gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G211gat), .ZN(new_n213_));
  INV_X1    g012(.A(G211gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G218gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT92), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n210_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(G204gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n209_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT21), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n205_), .A2(new_n208_), .A3(new_n211_), .A4(new_n209_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT26), .B(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228_));
  OR2_X1    g027(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT23), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n246_));
  INV_X1    g045(.A(new_n243_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n233_), .A2(new_n242_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n251_), .C1(KEYINPUT22), .C2(G176gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G190gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n229_), .A2(new_n258_), .A3(new_n230_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n259_), .B(new_n261_), .C1(new_n243_), .C2(new_n246_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n221_), .A2(new_n226_), .A3(new_n249_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT20), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT82), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n260_), .B1(new_n270_), .B2(new_n247_), .ZN(new_n271_));
  AND2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(new_n239_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n240_), .A2(KEYINPUT93), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n240_), .A2(KEYINPUT93), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n239_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT25), .B(G183gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n227_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n271_), .A2(new_n276_), .A3(new_n278_), .A4(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT22), .B(G169gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n272_), .B1(new_n282_), .B2(new_n235_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n244_), .B1(new_n270_), .B2(new_n243_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n210_), .A2(new_n219_), .A3(new_n216_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n219_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n226_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n203_), .B1(new_n265_), .B2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT20), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n249_), .A2(new_n263_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n290_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n203_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n213_), .A2(new_n215_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(KEYINPUT21), .B2(new_n223_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n218_), .A2(new_n220_), .B1(new_n225_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n293_), .A2(new_n297_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT27), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT100), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n238_), .A2(new_n241_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n284_), .A2(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n311_), .A2(new_n233_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n304_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n287_), .A2(new_n290_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n203_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT97), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n300_), .A2(new_n305_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(KEYINPUT97), .A3(new_n203_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n264_), .A2(new_n291_), .A3(KEYINPUT20), .A4(new_n301_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT98), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n298_), .B1(new_n312_), .B2(new_n304_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(KEYINPUT98), .A3(new_n301_), .A4(new_n291_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n317_), .A2(new_n319_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n297_), .B(KEYINPUT99), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n309_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n324_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT97), .B1(new_n318_), .B2(new_n203_), .ZN(new_n330_));
  AOI211_X1 g129(.A(new_n316_), .B(new_n301_), .C1(new_n300_), .C2(new_n305_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT100), .A3(new_n326_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n308_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n299_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n312_), .A2(KEYINPUT30), .ZN(new_n337_));
  INV_X1    g136(.A(G99gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n249_), .A2(new_n263_), .A3(KEYINPUT30), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT30), .B1(new_n249_), .B2(new_n263_), .ZN(new_n341_));
  OAI21_X1  g140(.A(G99gat), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G15gat), .B(G43gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G71gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n345_), .B(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n339_), .A2(new_n342_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT86), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n339_), .A2(new_n342_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n348_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n339_), .A2(new_n342_), .A3(new_n348_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT31), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n351_), .A2(new_n357_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT95), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT88), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(G155gat), .A3(G162gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n366_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OR3_X1    g176(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n371_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n368_), .A2(new_n370_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n385_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n366_), .ZN(new_n388_));
  OR3_X1    g187(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n379_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n365_), .B(new_n384_), .C1(new_n388_), .C2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(new_n362_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n362_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n368_), .A2(new_n370_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT1), .ZN(new_n397_));
  INV_X1    g196(.A(new_n366_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n368_), .A2(new_n370_), .A3(new_n385_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n391_), .A2(new_n379_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n376_), .A2(new_n378_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n400_), .A2(new_n401_), .B1(new_n402_), .B2(new_n371_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n395_), .B1(new_n403_), .B2(new_n365_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT4), .B1(new_n394_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n384_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n362_), .A2(KEYINPUT4), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n405_), .A2(new_n406_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n393_), .A2(new_n362_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n403_), .A2(new_n365_), .A3(new_n395_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT96), .B1(new_n418_), .B2(new_n412_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G57gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  AOI21_X1  g222(.A(new_n411_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n414_), .A2(new_n419_), .A3(new_n423_), .A4(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n414_), .A2(new_n419_), .A3(new_n425_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n423_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n363_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .A4(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n364_), .A2(new_n426_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(G78gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G106gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT28), .B1(new_n407_), .B2(KEYINPUT29), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n403_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n437_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n441_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT90), .ZN(new_n447_));
  INV_X1    g246(.A(new_n437_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n304_), .B1(KEYINPUT29), .B2(new_n407_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G22gat), .B(G50gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n445_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n297_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n313_), .A2(new_n203_), .A3(new_n314_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n301_), .B1(new_n323_), .B2(new_n291_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT94), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n307_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT27), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT94), .B(new_n457_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR4_X1   g265(.A1(new_n334_), .A2(new_n432_), .A3(new_n456_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n464_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n426_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n416_), .A2(new_n417_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n412_), .B1(new_n471_), .B2(KEYINPUT4), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n424_), .B1(new_n472_), .B2(new_n406_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n473_), .A2(KEYINPUT33), .A3(new_n423_), .A4(new_n419_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n423_), .B1(new_n471_), .B2(new_n411_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n409_), .A2(new_n410_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n418_), .B2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n468_), .A2(new_n470_), .A3(new_n474_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n332_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n293_), .A2(new_n479_), .A3(new_n306_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n423_), .B1(new_n473_), .B2(new_n419_), .ZN(new_n483_));
  AND4_X1   g282(.A1(new_n423_), .A2(new_n414_), .A3(new_n419_), .A4(new_n425_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n481_), .B(new_n482_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n454_), .A2(new_n455_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n308_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n325_), .A2(new_n309_), .A3(new_n327_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT100), .B1(new_n332_), .B2(new_n326_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n429_), .A2(new_n426_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n492_), .A2(new_n456_), .A3(new_n494_), .A4(new_n465_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n364_), .A2(new_n431_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n467_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT76), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G15gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(G22gat), .ZN(new_n507_));
  INV_X1    g306(.A(G22gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(G15gat), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n507_), .A2(new_n509_), .A3(KEYINPUT76), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G1gat), .A2(G8gat), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n511_), .A2(KEYINPUT77), .A3(KEYINPUT14), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT77), .B1(new_n511_), .B2(KEYINPUT14), .ZN(new_n513_));
  OAI22_X1  g312(.A1(new_n505_), .A2(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G1gat), .B(G8gat), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  OAI221_X1 g316(.A(new_n515_), .B1(new_n513_), .B2(new_n512_), .C1(new_n505_), .C2(new_n510_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G29gat), .B(G36gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT72), .ZN(new_n523_));
  INV_X1    g322(.A(G36gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G29gat), .ZN(new_n525_));
  INV_X1    g324(.A(G29gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G36gat), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n525_), .A2(new_n527_), .A3(KEYINPUT72), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n521_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n527_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(KEYINPUT72), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n520_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(KEYINPUT15), .A3(new_n534_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n519_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n517_), .A2(new_n535_), .A3(new_n518_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n517_), .A2(new_n535_), .A3(new_n518_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n535_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n546_), .A3(KEYINPUT78), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT78), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n539_), .A2(new_n548_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n502_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n502_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT79), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT79), .ZN(new_n554_));
  AND4_X1   g353(.A1(new_n554_), .A2(new_n547_), .A3(new_n549_), .A4(new_n502_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n556_), .A3(KEYINPUT80), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n498_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566_));
  INV_X1    g365(.A(G85gat), .ZN(new_n567_));
  INV_X1    g366(.A(G92gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n566_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n564_), .B(new_n566_), .C1(new_n570_), .C2(new_n569_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT10), .B(G99gat), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n436_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT6), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .A4(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT8), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n338_), .A3(new_n436_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n569_), .A2(new_n566_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n576_), .B(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n580_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n584_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(KEYINPUT8), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n578_), .B1(new_n585_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n535_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT73), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(KEYINPUT8), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n594_), .A2(new_n595_), .B1(new_n596_), .B2(new_n572_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n535_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n593_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT67), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n591_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT67), .B(new_n578_), .C1(new_n585_), .C2(new_n590_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n602_), .A2(new_n538_), .A3(new_n537_), .A4(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT34), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT35), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(KEYINPUT35), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT71), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n593_), .A2(new_n599_), .B1(new_n608_), .B2(new_n607_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n604_), .A3(new_n612_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT75), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n614_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n619_), .B(KEYINPUT36), .Z(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n563_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G57gat), .B(G64gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G71gat), .B(G78gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(KEYINPUT11), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(KEYINPUT11), .ZN(new_n630_));
  INV_X1    g429(.A(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n627_), .A2(KEYINPUT11), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n519_), .B(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n636_), .B(new_n637_), .Z(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT17), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n636_), .B(new_n637_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT17), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n624_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n616_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n612_), .B1(new_n615_), .B2(new_n604_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n614_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT37), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n626_), .A2(new_n649_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT66), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n597_), .A2(new_n657_), .A3(new_n634_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n578_), .B(new_n634_), .C1(new_n585_), .C2(new_n590_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT66), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n591_), .A2(new_n635_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT64), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n635_), .A2(KEYINPUT12), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n602_), .A2(new_n668_), .A3(new_n603_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT12), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n661_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n665_), .B1(new_n597_), .B2(new_n634_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n666_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(G120gat), .B(G148gat), .Z(new_n675_));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n677_), .B(new_n678_), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n666_), .A2(new_n673_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT69), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(KEYINPUT69), .A3(new_n682_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n680_), .A2(KEYINPUT69), .A3(new_n682_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT69), .B1(new_n680_), .B2(new_n682_), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n689_), .A2(new_n690_), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n656_), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n562_), .A2(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(G1gat), .A3(new_n494_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT38), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT38), .ZN(new_n696_));
  INV_X1    g495(.A(G1gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n691_), .A2(new_n688_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n547_), .A2(new_n549_), .A3(new_n502_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n555_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n701_), .A3(new_n649_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT101), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n429_), .B(new_n426_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n334_), .A2(new_n704_), .A3(new_n466_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n456_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n497_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n334_), .A2(new_n466_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n497_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n708_), .A2(new_n487_), .A3(new_n494_), .A4(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n623_), .A2(new_n625_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n703_), .A2(new_n494_), .A3(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n695_), .B(new_n696_), .C1(new_n697_), .C2(new_n715_), .ZN(G1324gat));
  INV_X1    g515(.A(G8gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n703_), .A2(new_n714_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n708_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT39), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n693_), .A2(G8gat), .A3(new_n708_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT102), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT40), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n722_), .A2(KEYINPUT40), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1325gat));
  AOI21_X1  g528(.A(new_n506_), .B1(new_n718_), .B2(new_n709_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT104), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n693_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n506_), .A3(new_n709_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n730_), .A2(new_n732_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n733_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT105), .ZN(G1326gat));
  AOI21_X1  g537(.A(new_n508_), .B1(new_n718_), .B2(new_n456_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT42), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n508_), .A3(new_n456_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1327gat));
  INV_X1    g541(.A(new_n698_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n743_), .A2(new_n649_), .A3(new_n713_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n562_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G29gat), .B1(new_n746_), .B2(new_n493_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n623_), .A2(new_n625_), .A3(new_n563_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT37), .B1(new_n653_), .B2(new_n654_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n498_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n752_));
  INV_X1    g551(.A(new_n750_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n711_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n743_), .A2(new_n557_), .A3(new_n649_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(KEYINPUT44), .A3(new_n756_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n494_), .A2(new_n526_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n747_), .B1(new_n761_), .B2(new_n762_), .ZN(G1328gat));
  NAND3_X1  g562(.A1(new_n746_), .A2(new_n524_), .A3(new_n719_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT45), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(new_n719_), .A3(new_n760_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G36gat), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(new_n767_), .A3(KEYINPUT46), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1329gat));
  NAND4_X1  g571(.A1(new_n759_), .A2(G43gat), .A3(new_n709_), .A4(new_n760_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n745_), .A2(new_n497_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(G43gat), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g575(.A1(new_n745_), .A2(G50gat), .A3(new_n487_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n761_), .A2(KEYINPUT106), .A3(new_n456_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G50gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT106), .B1(new_n761_), .B2(new_n456_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(G1331gat));
  NOR2_X1   g580(.A1(new_n498_), .A2(new_n712_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n743_), .A2(new_n561_), .A3(new_n649_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n494_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n656_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n698_), .A2(new_n701_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n711_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G57gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n493_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n791_), .ZN(G1332gat));
  INV_X1    g591(.A(G64gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n784_), .B2(new_n719_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT48), .Z(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n793_), .A3(new_n719_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1333gat));
  NOR2_X1   g596(.A1(new_n497_), .A2(G71gat), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT107), .Z(new_n799_));
  NAND2_X1  g598(.A1(new_n789_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n784_), .A2(new_n709_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G71gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G71gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1334gat));
  AOI21_X1  g606(.A(new_n434_), .B1(new_n784_), .B2(new_n456_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n789_), .A2(new_n434_), .A3(new_n456_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1335gat));
  NAND2_X1  g611(.A1(new_n644_), .A2(new_n648_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n711_), .A2(new_n813_), .A3(new_n712_), .A4(new_n788_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n815_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n493_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n818_), .A2(new_n567_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n819_), .A2(KEYINPUT111), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT111), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n698_), .A2(new_n701_), .A3(new_n649_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n494_), .A2(new_n567_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n820_), .A2(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(G1336gat));
  OAI21_X1  g625(.A(new_n719_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n708_), .A2(new_n568_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT112), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n827_), .A2(new_n568_), .B1(new_n824_), .B2(new_n829_), .ZN(G1337gat));
  OAI211_X1 g629(.A(new_n709_), .B(new_n574_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n824_), .A2(new_n709_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n338_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g633(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n752_), .B1(new_n711_), .B2(new_n753_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT43), .B(new_n750_), .C1(new_n707_), .C2(new_n710_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n456_), .B(new_n822_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G106gat), .B1(new_n839_), .B2(KEYINPUT113), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n824_), .B2(new_n456_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n836_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n824_), .A2(new_n841_), .A3(new_n456_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(KEYINPUT113), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(G106gat), .A4(new_n835_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n436_), .B(new_n456_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT53), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1339gat));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n669_), .A2(new_n671_), .A3(new_n660_), .A4(new_n658_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n665_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n669_), .A2(new_n671_), .A3(KEYINPUT55), .A4(new_n672_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n673_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n857_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n679_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(new_n679_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n682_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n685_), .A2(new_n686_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n539_), .A2(new_n541_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n540_), .B1(new_n867_), .B2(KEYINPUT115), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(KEYINPUT115), .B2(new_n867_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n540_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n502_), .A3(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(new_n551_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n865_), .A2(new_n701_), .B1(new_n866_), .B2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT116), .B(new_n854_), .C1(new_n873_), .C2(new_n712_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n860_), .A2(new_n679_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT56), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n860_), .A2(new_n861_), .A3(new_n679_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n701_), .A2(new_n876_), .A3(new_n682_), .A4(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n872_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n712_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT57), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n865_), .A2(KEYINPUT58), .A3(new_n872_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n876_), .A2(new_n682_), .A3(new_n872_), .A4(new_n877_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n753_), .A3(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n874_), .A2(new_n882_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n813_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n692_), .B2(new_n561_), .ZN(new_n891_));
  AND4_X1   g690(.A1(new_n890_), .A2(new_n787_), .A3(new_n698_), .A4(new_n561_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n719_), .A2(new_n456_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n493_), .A3(new_n709_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(KEYINPUT59), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n893_), .B1(new_n888_), .B2(new_n813_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n897_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n561_), .B1(new_n899_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(G113gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n895_), .A2(new_n898_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n557_), .A2(G113gat), .ZN(new_n906_));
  OAI22_X1  g705(.A1(new_n903_), .A2(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1340gat));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT117), .B(G120gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n899_), .A2(new_n902_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n743_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n901_), .A2(new_n897_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n909_), .A2(KEYINPUT60), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n698_), .A2(KEYINPUT60), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n915_), .B2(new_n909_), .ZN(new_n916_));
  AOI21_X1  g715(.A(KEYINPUT118), .B1(new_n912_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918_));
  INV_X1    g717(.A(new_n916_), .ZN(new_n919_));
  NOR4_X1   g718(.A1(new_n901_), .A2(new_n918_), .A3(new_n897_), .A4(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n908_), .B1(new_n911_), .B2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n698_), .B1(new_n899_), .B2(new_n902_), .ZN(new_n923_));
  OAI221_X1 g722(.A(KEYINPUT119), .B1(new_n917_), .B2(new_n920_), .C1(new_n923_), .C2(new_n909_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1341gat));
  INV_X1    g724(.A(G127gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n905_), .B2(new_n813_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n813_), .A2(new_n926_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n930_), .B1(new_n910_), .B2(new_n931_), .ZN(G1342gat));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933_));
  INV_X1    g732(.A(G134gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n910_), .B2(new_n753_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n712_), .A2(new_n934_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n905_), .A2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n933_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n750_), .B1(new_n899_), .B2(new_n902_), .ZN(new_n939_));
  OAI221_X1 g738(.A(KEYINPUT121), .B1(new_n905_), .B2(new_n936_), .C1(new_n939_), .C2(new_n934_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1343gat));
  NOR3_X1   g740(.A1(new_n709_), .A2(new_n494_), .A3(new_n487_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n895_), .A2(new_n708_), .A3(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n557_), .ZN(new_n944_));
  XOR2_X1   g743(.A(new_n944_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g744(.A1(new_n943_), .A2(new_n698_), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n946_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g746(.A1(new_n943_), .A2(new_n813_), .ZN(new_n948_));
  XOR2_X1   g747(.A(KEYINPUT61), .B(G155gat), .Z(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1346gat));
  OAI21_X1  g749(.A(G162gat), .B1(new_n943_), .B2(new_n750_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n713_), .A2(G162gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n943_), .B2(new_n952_), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n901_), .A2(new_n708_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n432_), .A2(new_n456_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  OAI21_X1  g755(.A(G169gat), .B1(new_n956_), .B2(new_n557_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n954_), .A2(new_n282_), .A3(new_n701_), .A4(new_n955_), .ZN(new_n960_));
  OAI211_X1 g759(.A(KEYINPUT62), .B(G169gat), .C1(new_n956_), .C2(new_n557_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(G1348gat));
  NOR2_X1   g761(.A1(new_n956_), .A2(new_n698_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n235_), .A2(KEYINPUT122), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  XOR2_X1   g764(.A(KEYINPUT122), .B(G176gat), .Z(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n963_), .B2(new_n966_), .ZN(G1349gat));
  NOR2_X1   g766(.A1(new_n956_), .A2(new_n813_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n229_), .A2(new_n230_), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n968_), .B(new_n279_), .C1(KEYINPUT123), .C2(new_n969_), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n229_), .A2(KEYINPUT123), .A3(new_n230_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n968_), .B2(new_n971_), .ZN(G1350gat));
  OAI21_X1  g771(.A(G190gat), .B1(new_n956_), .B2(new_n750_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n712_), .A2(new_n227_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n956_), .B2(new_n974_), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n709_), .A2(new_n704_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n954_), .A2(new_n976_), .ZN(new_n977_));
  INV_X1    g776(.A(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978_), .B2(new_n701_), .ZN(new_n979_));
  NAND4_X1  g778(.A1(new_n954_), .A2(G197gat), .A3(new_n701_), .A4(new_n976_), .ZN(new_n980_));
  AND2_X1   g779(.A1(new_n980_), .A2(KEYINPUT124), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n980_), .A2(KEYINPUT124), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n979_), .A2(new_n981_), .A3(new_n982_), .ZN(G1352gat));
  OAI21_X1  g782(.A(new_n743_), .B1(KEYINPUT125), .B2(new_n204_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n977_), .A2(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n204_), .A2(KEYINPUT125), .ZN(new_n986_));
  XOR2_X1   g785(.A(new_n986_), .B(KEYINPUT126), .Z(new_n987_));
  XNOR2_X1  g786(.A(new_n985_), .B(new_n987_), .ZN(G1353gat));
  AOI211_X1 g787(.A(KEYINPUT63), .B(G211gat), .C1(new_n978_), .C2(new_n649_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(KEYINPUT63), .B(G211gat), .ZN(new_n990_));
  NOR3_X1   g789(.A1(new_n977_), .A2(new_n813_), .A3(new_n990_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n989_), .A2(new_n991_), .ZN(G1354gat));
  NOR3_X1   g791(.A1(new_n977_), .A2(new_n212_), .A3(new_n750_), .ZN(new_n993_));
  NOR3_X1   g792(.A1(new_n977_), .A2(KEYINPUT127), .A3(new_n713_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(new_n994_), .A2(G218gat), .ZN(new_n995_));
  OAI21_X1  g794(.A(KEYINPUT127), .B1(new_n977_), .B2(new_n713_), .ZN(new_n996_));
  AOI21_X1  g795(.A(new_n993_), .B1(new_n995_), .B2(new_n996_), .ZN(G1355gat));
endmodule


