//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT30), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT31), .ZN(new_n206_));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207_));
  XOR2_X1   g006(.A(G113gat), .B(G120gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT22), .B(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n211_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT82), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n212_), .A2(KEYINPUT81), .A3(new_n213_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n216_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n220_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n211_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(G183gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n237_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT26), .B(G190gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT80), .B1(new_n237_), .B2(KEYINPUT25), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n232_), .B(new_n233_), .C1(new_n236_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n227_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT83), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n227_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  INV_X1    g048(.A(G43gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n247_), .A2(new_n251_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n209_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n209_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n206_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n206_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n259_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT84), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G1gat), .B(G29gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G85gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT0), .B(G57gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT95), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G225gat), .A2(G233gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT86), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n273_), .A2(new_n275_), .B1(new_n276_), .B2(KEYINPUT85), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n271_), .B1(new_n274_), .B2(new_n272_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(KEYINPUT2), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n280_), .A2(new_n274_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n276_), .A2(KEYINPUT85), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n277_), .A2(new_n278_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n281_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n274_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n286_), .A2(KEYINPUT1), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(KEYINPUT1), .B2(new_n286_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n209_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n295_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n209_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT93), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT93), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n299_), .A2(new_n305_), .A3(KEYINPUT4), .A4(new_n301_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n297_), .A2(new_n303_), .A3(new_n298_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT94), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n270_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n302_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n270_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n267_), .B(new_n269_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT95), .B1(new_n316_), .B2(new_n268_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n314_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n308_), .B(KEYINPUT94), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n322_), .B2(new_n270_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(new_n267_), .A3(new_n269_), .A4(new_n317_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n307_), .A2(new_n270_), .A3(new_n310_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n267_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT25), .B(G183gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n239_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n233_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n222_), .A2(new_n231_), .A3(new_n224_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT92), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n222_), .A2(new_n338_), .A3(new_n231_), .A4(new_n224_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n228_), .A2(new_n223_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G197gat), .B(G204gat), .Z(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n346_));
  XOR2_X1   g145(.A(G211gat), .B(G218gat), .Z(new_n347_));
  OAI22_X1  g146(.A1(new_n346_), .A2(new_n347_), .B1(KEYINPUT21), .B2(new_n345_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n344_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT19), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n344_), .B2(new_n350_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n244_), .A2(new_n246_), .A3(new_n352_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n332_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n355_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n353_), .A2(new_n355_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n351_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n367_), .A3(new_n331_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n327_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n319_), .A2(new_n324_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n353_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n350_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT97), .B1(new_n372_), .B2(new_n358_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n374_), .B(KEYINPUT20), .C1(new_n344_), .C2(new_n350_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(KEYINPUT98), .A3(new_n355_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n359_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n376_), .A2(new_n355_), .B1(new_n379_), .B2(KEYINPUT98), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT32), .B(new_n331_), .C1(new_n378_), .C2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n267_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n267_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n383_), .B(new_n320_), .C1(new_n322_), .C2(new_n270_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n364_), .A2(new_n367_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n370_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT89), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n392_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G22gat), .B(G50gat), .Z(new_n395_));
  OR3_X1    g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n352_), .B1(G228gat), .B2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n300_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G78gat), .B(G106gat), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n404_));
  OAI21_X1  g203(.A(new_n350_), .B1(new_n300_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(G228gat), .A3(G233gat), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n401_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n403_), .B1(new_n401_), .B2(new_n406_), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n398_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n398_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n389_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n368_), .A2(KEYINPUT27), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n353_), .B1(new_n351_), .B2(KEYINPUT97), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n357_), .B1(new_n415_), .B2(new_n375_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n379_), .A2(KEYINPUT98), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n377_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n418_), .B2(new_n332_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT27), .B1(new_n368_), .B2(new_n362_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n385_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n411_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n263_), .B1(new_n413_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT99), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n420_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n380_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n331_), .B1(new_n428_), .B2(new_n377_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n427_), .B(KEYINPUT99), .C1(new_n429_), .C2(new_n414_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n385_), .A2(new_n261_), .A3(new_n258_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n412_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT100), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n411_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT100), .A3(new_n432_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n424_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G1gat), .B(G8gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G22gat), .ZN(new_n442_));
  INV_X1    g241(.A(G1gat), .ZN(new_n443_));
  INV_X1    g242(.A(G8gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT14), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n441_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G29gat), .B(G36gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G43gat), .B(G50gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G43gat), .B(G50gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n448_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n441_), .B(new_n446_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n452_), .A2(KEYINPUT15), .A3(new_n454_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT15), .B1(new_n452_), .B2(new_n454_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n448_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n458_), .B2(new_n455_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n460_), .A2(new_n462_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G113gat), .B(G141gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G169gat), .B(G197gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  OR2_X1    g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n469_), .A2(KEYINPUT78), .A3(new_n472_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT78), .B1(new_n469_), .B2(new_n472_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n438_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G231gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(G71gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT64), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT64), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(G71gat), .ZN(new_n483_));
  INV_X1    g282(.A(G78gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(KEYINPUT11), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT64), .B(G71gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(new_n484_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT65), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(new_n483_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G78gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT11), .ZN(new_n493_));
  INV_X1    g292(.A(G57gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(G64gat), .ZN(new_n495_));
  INV_X1    g294(.A(G64gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(G57gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n493_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n492_), .A2(new_n498_), .A3(new_n499_), .A4(new_n485_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(G57gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(G64gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(new_n493_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n490_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n490_), .B2(new_n500_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n479_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n479_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT76), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n508_), .A2(KEYINPUT76), .A3(new_n509_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n511_), .A2(new_n458_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G127gat), .B(G155gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(G183gat), .B(G211gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n458_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n514_), .A2(KEYINPUT17), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n519_), .B(KEYINPUT17), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n513_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT6), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n530_));
  OR2_X1    g329(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G85gat), .ZN(new_n535_));
  INV_X1    g334(.A(G92gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(KEYINPUT9), .A3(new_n529_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n528_), .A2(new_n530_), .A3(new_n534_), .A4(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n537_), .A2(new_n529_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n527_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544_));
  INV_X1    g343(.A(G99gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n532_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n541_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT8), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n542_), .B1(G99gat), .B2(G106gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n527_), .A2(KEYINPUT6), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n547_), .B(new_n546_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT8), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n541_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n540_), .B1(new_n550_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT34), .Z(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n556_), .A2(new_n455_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n455_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n463_), .ZN(new_n563_));
  OAI221_X1 g362(.A(new_n560_), .B1(new_n563_), .B2(new_n556_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n556_), .B2(new_n563_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n555_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n554_), .B1(new_n553_), .B2(new_n541_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n539_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n466_), .A3(KEYINPUT70), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n560_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n558_), .A2(new_n559_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(KEYINPUT71), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT71), .B1(new_n576_), .B2(new_n577_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n564_), .B(new_n569_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n564_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n567_), .B(KEYINPUT36), .Z(new_n584_));
  AND3_X1   g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n583_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n580_), .B(new_n581_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n582_), .A2(new_n584_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n580_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT37), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n526_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT66), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n574_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n504_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n493_), .A2(new_n503_), .B1(new_n488_), .B2(new_n484_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n499_), .B1(new_n595_), .B2(new_n492_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n500_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n490_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n556_), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n600_), .A3(KEYINPUT12), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n574_), .B(new_n602_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n592_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  AOI211_X1 g406(.A(KEYINPUT66), .B(new_n607_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n605_), .B1(new_n593_), .B2(new_n600_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n606_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT67), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT68), .B1(new_n610_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n604_), .A2(new_n605_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT66), .ZN(new_n619_));
  INV_X1    g418(.A(new_n609_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n607_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n592_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .A4(new_n614_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT68), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n615_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n617_), .A2(new_n623_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT13), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n617_), .A2(KEYINPUT13), .A3(new_n623_), .A4(new_n626_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n478_), .A2(new_n591_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n443_), .A3(new_n385_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT104), .Z(new_n636_));
  INV_X1    g435(.A(new_n526_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n631_), .A2(new_n476_), .A3(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT102), .Z(new_n639_));
  OAI21_X1  g438(.A(new_n580_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT103), .Z(new_n641_));
  NOR2_X1   g440(.A1(new_n438_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n422_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n636_), .B(new_n644_), .C1(new_n634_), .C2(new_n633_), .ZN(G1324gat));
  INV_X1    g444(.A(new_n431_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n632_), .A2(new_n444_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G8gat), .B1(new_n643_), .B2(new_n431_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT39), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT39), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n651_), .B(new_n653_), .ZN(G1325gat));
  NAND3_X1  g453(.A1(new_n639_), .A2(new_n263_), .A3(new_n642_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G15gat), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT106), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT106), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(KEYINPUT41), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n632_), .A2(new_n203_), .A3(new_n263_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(new_n657_), .B2(new_n658_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n643_), .B2(new_n412_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n412_), .A2(G22gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT107), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n632_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n631_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n670_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n478_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n385_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n631_), .A2(new_n476_), .A3(new_n526_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n587_), .A2(new_n590_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n438_), .A2(KEYINPUT43), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(new_n263_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n423_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n411_), .B1(new_n370_), .B2(new_n388_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AND4_X1   g481(.A1(KEYINPUT100), .A2(new_n431_), .A3(new_n412_), .A4(new_n432_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT100), .B1(new_n436_), .B2(new_n432_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n676_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n678_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n675_), .B1(new_n677_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n438_), .B2(new_n676_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n685_), .A2(new_n678_), .A3(new_n686_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n674_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n690_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(KEYINPUT44), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n385_), .A2(G29gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n673_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n431_), .B1(new_n693_), .B2(KEYINPUT44), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n696_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n672_), .A2(new_n705_), .A3(new_n646_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n703_), .B(new_n704_), .C1(new_n707_), .C2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n695_), .B1(new_n693_), .B2(KEYINPUT108), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n688_), .A2(new_n689_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n706_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n715_), .A2(new_n701_), .A3(new_n716_), .A4(new_n702_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n711_), .A2(new_n717_), .ZN(G1329gat));
  NAND4_X1  g517(.A1(new_n696_), .A2(G43gat), .A3(new_n262_), .A4(new_n697_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n672_), .A2(new_n263_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n250_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n719_), .A2(KEYINPUT47), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT47), .B1(new_n719_), .B2(new_n721_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n672_), .B2(new_n411_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n411_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n698_), .B2(new_n726_), .ZN(G1331gat));
  NAND4_X1  g526(.A1(new_n642_), .A2(new_n477_), .A3(new_n637_), .A4(new_n670_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n422_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n670_), .A2(new_n477_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n438_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n591_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n385_), .A2(new_n494_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1332gat));
  OAI21_X1  g533(.A(G64gat), .B1(new_n728_), .B2(new_n431_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT48), .ZN(new_n736_));
  INV_X1    g535(.A(new_n732_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n496_), .A3(new_n646_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n728_), .B2(new_n679_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT49), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n263_), .A2(new_n480_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT110), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n732_), .B2(new_n743_), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n728_), .B2(new_n412_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n484_), .A3(new_n411_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1335gat));
  NAND3_X1  g547(.A1(new_n670_), .A2(new_n477_), .A3(new_n526_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n422_), .ZN(new_n752_));
  NOR4_X1   g551(.A1(new_n438_), .A2(new_n730_), .A3(new_n640_), .A4(new_n637_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n535_), .A3(new_n385_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1336gat));
  OAI21_X1  g554(.A(G92gat), .B1(new_n751_), .B2(new_n431_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n536_), .A3(new_n646_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1337gat));
  NAND4_X1  g557(.A1(new_n753_), .A2(new_n262_), .A3(new_n531_), .A4(new_n533_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(KEYINPUT111), .B2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n545_), .B1(new_n750_), .B2(new_n263_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(KEYINPUT111), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n763_), .B(new_n764_), .Z(G1338gat));
  NAND3_X1  g564(.A1(new_n753_), .A2(new_n532_), .A3(new_n411_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n411_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G106gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT52), .B(new_n532_), .C1(new_n750_), .C2(new_n411_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1339gat));
  NAND3_X1  g572(.A1(new_n436_), .A2(new_n262_), .A3(new_n385_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT117), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n591_), .A2(new_n477_), .A3(new_n629_), .A4(new_n630_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT113), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT113), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n631_), .A2(new_n781_), .A3(new_n477_), .A4(new_n591_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n777_), .A2(KEYINPUT113), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT54), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n780_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT114), .B1(new_n623_), .B2(new_n476_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n623_), .A2(new_n476_), .A3(KEYINPUT114), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n619_), .A2(new_n622_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n601_), .A2(new_n607_), .A3(new_n603_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(KEYINPUT55), .B2(new_n621_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n615_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n796_), .B(new_n616_), .C1(new_n790_), .C2(new_n793_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n787_), .B(new_n788_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n474_), .A2(new_n475_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n467_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n472_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n627_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT57), .B1(new_n804_), .B2(new_n640_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  INV_X1    g605(.A(new_n640_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n806_), .B(new_n807_), .C1(new_n798_), .C2(new_n803_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n789_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n606_), .A2(new_n608_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n791_), .B1(new_n618_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT56), .B(new_n615_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT116), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n794_), .A2(new_n816_), .A3(KEYINPUT56), .A4(new_n615_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n606_), .A2(new_n608_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n813_), .B1(new_n818_), .B2(new_n789_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n796_), .B1(new_n819_), .B2(new_n616_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n802_), .A2(new_n623_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT58), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n676_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n821_), .A2(KEYINPUT58), .A3(new_n822_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n637_), .B1(new_n809_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n775_), .B1(new_n785_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n476_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  INV_X1    g632(.A(new_n775_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n782_), .A2(KEYINPUT54), .A3(new_n783_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT54), .B1(new_n782_), .B2(new_n783_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n788_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n786_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n820_), .A2(new_n814_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n839_), .A2(new_n840_), .B1(new_n627_), .B2(new_n802_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n806_), .B1(new_n841_), .B2(new_n807_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n804_), .A2(KEYINPUT57), .A3(new_n640_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n825_), .A2(new_n823_), .A3(new_n676_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n526_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n833_), .B(new_n834_), .C1(new_n837_), .C2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n784_), .A3(new_n780_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT59), .B1(new_n848_), .B2(new_n775_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n832_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n829_), .A2(new_n833_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(KEYINPUT59), .A3(new_n775_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(KEYINPUT118), .A3(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(G113gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n477_), .A2(new_n855_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT120), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n831_), .B1(new_n854_), .B2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n631_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n830_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n631_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n859_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n526_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n850_), .A2(new_n853_), .A3(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n829_), .B2(new_n526_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n866_), .A2(KEYINPUT121), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT121), .B1(new_n866_), .B2(new_n867_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1342gat));
  NAND3_X1  g669(.A1(new_n850_), .A2(new_n686_), .A3(new_n853_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G134gat), .ZN(new_n872_));
  INV_X1    g671(.A(new_n641_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n873_), .A2(G134gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n829_), .B2(new_n874_), .ZN(G1343gat));
  NOR2_X1   g674(.A1(new_n263_), .A2(new_n412_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n848_), .A2(new_n385_), .A3(new_n431_), .A4(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n477_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT122), .B(G141gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1344gat));
  NOR2_X1   g679(.A1(new_n877_), .A2(new_n631_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g681(.A1(new_n877_), .A2(new_n526_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT61), .B(G155gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  OAI21_X1  g684(.A(G162gat), .B1(new_n877_), .B2(new_n676_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n873_), .A2(G162gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n877_), .B2(new_n887_), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n785_), .A2(new_n828_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n431_), .A2(new_n385_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n263_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n889_), .A2(new_n411_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n476_), .A2(new_n212_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT124), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n891_), .A2(new_n477_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT123), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n848_), .A2(new_n412_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n895_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT125), .ZN(G1348gat));
  NAND2_X1  g702(.A1(new_n892_), .A2(new_n670_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT126), .B(G176gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1349gat));
  NAND2_X1  g705(.A1(new_n892_), .A2(new_n637_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n333_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n237_), .B2(new_n907_), .ZN(G1350gat));
  INV_X1    g708(.A(new_n892_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G190gat), .B1(new_n910_), .B2(new_n676_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n892_), .A2(new_n239_), .A3(new_n641_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1351gat));
  NAND2_X1  g712(.A1(new_n876_), .A2(new_n890_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n889_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n476_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n670_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n637_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  NAND2_X1  g723(.A1(new_n915_), .A2(new_n686_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n873_), .A2(G218gat), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n925_), .A2(G218gat), .B1(new_n915_), .B2(new_n926_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


