//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_;
  XOR2_X1   g000(.A(G120gat), .B(G148gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G176gat), .B(G204gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n209_));
  OR3_X1    g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT11), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n207_), .B(KEYINPUT67), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT11), .ZN(new_n212_));
  XOR2_X1   g011(.A(G71gat), .B(G78gat), .Z(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n213_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(KEYINPUT11), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT12), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n223_), .B(new_n224_), .C1(new_n225_), .C2(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n222_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(KEYINPUT7), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT65), .A4(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT6), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT6), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(G99gat), .A3(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n221_), .B1(new_n235_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n239_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n229_), .A2(new_n233_), .A3(new_n246_), .A4(new_n234_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT8), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n221_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(KEYINPUT70), .A3(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT10), .B(G99gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n224_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n254_));
  INV_X1    g053(.A(G85gat), .ZN(new_n255_));
  INV_X1    g054(.A(G92gat), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n255_), .A2(new_n256_), .A3(KEYINPUT9), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n253_), .A2(new_n254_), .A3(new_n246_), .A4(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n244_), .A2(KEYINPUT8), .B1(new_n247_), .B2(new_n249_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT70), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n220_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n258_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n260_), .B2(KEYINPUT70), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n246_), .A2(KEYINPUT66), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n233_), .A2(new_n234_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n229_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n248_), .B1(new_n270_), .B2(new_n221_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n250_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n265_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n264_), .A2(KEYINPUT71), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n219_), .B1(new_n262_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n258_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT12), .B1(new_n218_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G230gat), .ZN(new_n278_));
  INV_X1    g077(.A(G233gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n260_), .A2(new_n263_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(new_n217_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n275_), .A2(new_n277_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n280_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT69), .B1(new_n281_), .B2(new_n217_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n218_), .A2(new_n276_), .A3(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n218_), .A2(new_n276_), .A3(KEYINPUT68), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n281_), .B2(new_n217_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n285_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n206_), .B1(new_n284_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n289_), .A2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n280_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n219_), .ZN(new_n299_));
  AND4_X1   g098(.A1(KEYINPUT71), .A2(new_n273_), .A3(new_n258_), .A4(new_n251_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT71), .B1(new_n264_), .B2(new_n273_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n277_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n282_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n206_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n298_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n295_), .A2(new_n296_), .A3(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(KEYINPUT73), .B(new_n206_), .C1(new_n284_), .C2(new_n294_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(KEYINPUT13), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(KEYINPUT13), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G29gat), .B(G36gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT75), .ZN(new_n314_));
  XOR2_X1   g113(.A(G43gat), .B(G50gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT15), .ZN(new_n317_));
  XOR2_X1   g116(.A(G15gat), .B(G22gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT78), .B(G1gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G8gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n320_), .B2(KEYINPUT14), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT79), .Z(new_n322_));
  XOR2_X1   g121(.A(G1gat), .B(G8gat), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(KEYINPUT79), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n323_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n327_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n316_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G229gat), .A2(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G113gat), .B(G141gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT83), .ZN(new_n335_));
  XOR2_X1   g134(.A(G169gat), .B(G197gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339_));
  INV_X1    g138(.A(new_n316_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n325_), .A2(new_n327_), .A3(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n330_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n339_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n333_), .B(new_n338_), .C1(new_n344_), .C2(new_n332_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n332_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n332_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n337_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n312_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(KEYINPUT21), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(KEYINPUT21), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G169gat), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n366_), .A2(KEYINPUT89), .A3(KEYINPUT22), .ZN(new_n367_));
  INV_X1    g166(.A(G176gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT22), .B1(new_n366_), .B2(KEYINPUT89), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT84), .B(G183gat), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(KEYINPUT23), .Z(new_n375_));
  OAI221_X1 g174(.A(new_n370_), .B1(new_n366_), .B2(new_n368_), .C1(new_n373_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n366_), .A2(new_n368_), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n380_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n371_), .A2(KEYINPUT25), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT85), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT26), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(G183gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT86), .B1(new_n386_), .B2(KEYINPUT25), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(G183gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(G190gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n387_), .B(new_n390_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  AOI211_X1 g192(.A(new_n385_), .B(new_n393_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n383_), .A2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n379_), .B(new_n381_), .C1(new_n395_), .C2(KEYINPUT88), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n383_), .A2(new_n394_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n365_), .B(new_n376_), .C1(new_n396_), .C2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G169gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n380_), .B1(new_n401_), .B2(new_n368_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n375_), .B2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT102), .Z(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT25), .B(G183gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT100), .ZN(new_n407_));
  INV_X1    g206(.A(new_n385_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n408_), .A2(new_n392_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n381_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT101), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n405_), .B1(new_n412_), .B2(new_n379_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n400_), .B(KEYINPUT20), .C1(new_n413_), .C2(new_n365_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT19), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n376_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n364_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT20), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(new_n379_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n365_), .A2(new_n404_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n418_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n358_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(new_n416_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n413_), .A2(new_n365_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n420_), .A2(new_n428_), .A3(KEYINPUT20), .A4(new_n418_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT0), .ZN(new_n432_));
  INV_X1    g231(.A(G57gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(new_n255_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT104), .ZN(new_n438_));
  INV_X1    g237(.A(G155gat), .ZN(new_n439_));
  INV_X1    g238(.A(G162gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n440_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G141gat), .A2(G148gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n443_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(new_n441_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n445_), .A2(new_n446_), .B1(KEYINPUT2), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G141gat), .A2(G148gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT94), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(KEYINPUT95), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT3), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT96), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G113gat), .B(G120gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT91), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G127gat), .B(G134gat), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(KEYINPUT92), .A3(new_n463_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n438_), .B1(new_n460_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n459_), .A2(KEYINPUT104), .A3(new_n469_), .A4(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n467_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n460_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT4), .A4(new_n474_), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n460_), .A2(new_n470_), .A3(KEYINPUT4), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n437_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n437_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n474_), .A2(new_n472_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n471_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n436_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n436_), .ZN(new_n483_));
  OAI221_X1 g282(.A(new_n426_), .B1(new_n430_), .B2(new_n358_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(KEYINPUT105), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT33), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n427_), .A2(new_n429_), .A3(new_n356_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT103), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n437_), .B1(new_n479_), .B2(new_n471_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n435_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT103), .ZN(new_n493_));
  INV_X1    g292(.A(new_n356_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n430_), .B2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n489_), .B(new_n492_), .C1(new_n495_), .C2(new_n488_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n484_), .B1(new_n486_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n470_), .B(KEYINPUT31), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n419_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504_));
  INV_X1    g303(.A(G43gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(G15gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n506_), .B(new_n509_), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n419_), .A2(new_n502_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n503_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n499_), .A2(new_n498_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n503_), .B2(new_n511_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n501_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n501_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n512_), .A3(new_n513_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G228gat), .A2(G233gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT97), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT98), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n364_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n524_), .B(new_n527_), .C1(new_n460_), .C2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n523_), .B1(new_n530_), .B2(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT99), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(KEYINPUT99), .A3(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(new_n539_), .A3(new_n531_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n460_), .A2(new_n541_), .A3(new_n528_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT28), .B1(new_n459_), .B2(KEYINPUT29), .ZN(new_n543_));
  XOR2_X1   g342(.A(G22gat), .B(G50gat), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n542_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n540_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n538_), .B(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n521_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n497_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n520_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n546_), .A2(new_n547_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n538_), .A2(new_n553_), .A3(new_n540_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n536_), .A2(new_n548_), .A3(new_n537_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n494_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n559_), .A2(KEYINPUT27), .A3(new_n487_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n489_), .B1(new_n495_), .B2(new_n488_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT27), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n482_), .A2(new_n483_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n551_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n352_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n217_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n329_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n571_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n571_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT80), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT80), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT81), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  OAI22_X1  g385(.A1(new_n276_), .A2(new_n340_), .B1(KEYINPUT35), .B2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n316_), .B(KEYINPUT15), .Z(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n274_), .B2(new_n262_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n590_));
  AOI211_X1 g389(.A(new_n587_), .B(new_n589_), .C1(KEYINPUT76), .C2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n589_), .B2(KEYINPUT76), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(new_n587_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n591_), .A2(new_n594_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n598_), .B(new_n600_), .C1(new_n591_), .C2(new_n594_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n603_));
  NOR2_X1   g402(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n583_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n568_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n564_), .A2(KEYINPUT106), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n564_), .A2(KEYINPUT106), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n610_), .A2(new_n319_), .A3(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT38), .Z(new_n616_));
  INV_X1    g415(.A(KEYINPUT107), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n352_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n602_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n551_), .B2(new_n566_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n582_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n565_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n622_), .ZN(G1324gat));
  OAI21_X1  g422(.A(G8gat), .B1(new_n621_), .B2(new_n563_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT39), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n610_), .A2(G8gat), .A3(new_n563_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(G1325gat));
  NOR3_X1   g428(.A1(new_n610_), .A2(G15gat), .A3(new_n520_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT108), .Z(new_n631_));
  NOR2_X1   g430(.A1(new_n621_), .A2(new_n520_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n632_), .A2(KEYINPUT41), .A3(new_n508_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT41), .B1(new_n632_), .B2(new_n508_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n633_), .A3(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n621_), .B2(new_n556_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT42), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n556_), .A2(G22gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n610_), .B2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n583_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n602_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n568_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n564_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n567_), .A2(new_n608_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n608_), .B2(KEYINPUT109), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n567_), .B(new_n608_), .C1(KEYINPUT109), .C2(new_n645_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n640_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n618_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(G29gat), .A3(new_n613_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n618_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n643_), .B1(new_n651_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(G36gat), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n563_), .A2(KEYINPUT111), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n563_), .A2(KEYINPUT111), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n642_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n563_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n654_), .A2(new_n663_), .A3(new_n650_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(new_n656_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1329gat));
  NOR2_X1   g466(.A1(new_n520_), .A2(new_n505_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n654_), .A2(new_n650_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT113), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT113), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n654_), .A2(new_n671_), .A3(new_n650_), .A4(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n642_), .A2(new_n521_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n505_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n642_), .B2(new_n549_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n650_), .A2(G50gat), .A3(new_n549_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n654_), .ZN(G1331gat));
  INV_X1    g482(.A(new_n312_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n350_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(new_n620_), .A3(new_n640_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(G57gat), .A3(new_n564_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT114), .Z(new_n688_));
  AND2_X1   g487(.A1(new_n685_), .A2(new_n567_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n609_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n433_), .B1(new_n690_), .B2(new_n614_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT115), .Z(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n686_), .B2(new_n659_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT48), .Z(new_n696_));
  INV_X1    g495(.A(new_n690_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n694_), .A3(new_n659_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n686_), .B2(new_n521_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT49), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n700_), .A3(new_n521_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT116), .ZN(G1334gat));
  INV_X1    g504(.A(G78gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n686_), .B2(new_n549_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT50), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n697_), .A2(new_n706_), .A3(new_n549_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1335gat));
  AND2_X1   g509(.A1(new_n649_), .A2(new_n685_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G85gat), .B1(new_n712_), .B2(new_n565_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n689_), .A2(new_n641_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n255_), .A3(new_n613_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1336gat));
  INV_X1    g516(.A(new_n659_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G92gat), .B1(new_n712_), .B2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n256_), .A3(new_n663_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1337gat));
  AOI21_X1  g520(.A(new_n223_), .B1(new_n711_), .B2(new_n521_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n521_), .A2(new_n252_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n715_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g524(.A1(new_n715_), .A2(new_n224_), .A3(new_n549_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n711_), .A2(new_n549_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G106gat), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT52), .B(new_n224_), .C1(new_n711_), .C2(new_n549_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(G1339gat));
  INV_X1    g532(.A(new_n582_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n333_), .B1(new_n344_), .B2(new_n332_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n331_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n337_), .B1(new_n736_), .B2(new_n347_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n344_), .A2(new_n332_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n735_), .A2(new_n337_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n307_), .A2(new_n739_), .A3(new_n308_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n302_), .A2(new_n303_), .A3(new_n293_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n280_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n304_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n302_), .A2(KEYINPUT55), .A3(new_n303_), .A4(new_n282_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n206_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n350_), .A2(new_n306_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT118), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n747_), .B2(new_n206_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n741_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n602_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n750_), .B1(new_n754_), .B2(KEYINPUT56), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n744_), .A2(new_n304_), .B1(new_n742_), .B2(new_n280_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n305_), .B1(new_n761_), .B2(new_n746_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n762_), .B2(new_n753_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n740_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT57), .B1(new_n764_), .B2(new_n619_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n758_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n747_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n206_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n748_), .A2(new_n760_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n739_), .A2(new_n306_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT58), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(KEYINPUT58), .A3(new_n773_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n608_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n777_), .A3(KEYINPUT120), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT120), .B1(new_n766_), .B2(new_n777_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n734_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n312_), .A2(new_n350_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n609_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n609_), .B2(new_n782_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n781_), .A2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n614_), .A2(new_n663_), .A3(new_n557_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n757_), .B1(new_n756_), .B2(new_n602_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n764_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n776_), .A2(new_n608_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n792_), .A2(new_n793_), .B1(new_n774_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n583_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n787_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n789_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n791_), .A2(new_n350_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G113gat), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT121), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n790_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n788_), .A2(KEYINPUT121), .A3(new_n789_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n351_), .A2(G113gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n801_), .A2(new_n806_), .ZN(G1340gat));
  NAND3_X1  g606(.A1(new_n791_), .A2(new_n312_), .A3(new_n799_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT122), .B(G120gat), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT60), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n312_), .A2(new_n812_), .A3(new_n809_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n812_), .B2(new_n809_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n803_), .A2(new_n804_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(G1341gat));
  AND2_X1   g615(.A1(new_n791_), .A2(new_n799_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n582_), .A2(G127gat), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT123), .Z(new_n819_));
  NAND3_X1  g618(.A1(new_n803_), .A2(new_n640_), .A3(new_n804_), .ZN(new_n820_));
  INV_X1    g619(.A(G127gat), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n817_), .A2(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(G1342gat));
  NAND3_X1  g621(.A1(new_n791_), .A2(new_n608_), .A3(new_n799_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G134gat), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n602_), .A2(G134gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n803_), .A2(new_n804_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1343gat));
  AOI21_X1  g626(.A(new_n552_), .B1(new_n781_), .B2(new_n787_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n613_), .A3(new_n718_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n350_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n312_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g633(.A1(new_n829_), .A2(new_n583_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT61), .B(G155gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  INV_X1    g636(.A(new_n608_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G162gat), .B1(new_n829_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n619_), .A2(new_n440_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n829_), .B2(new_n840_), .ZN(G1347gat));
  NOR3_X1   g640(.A1(new_n718_), .A2(new_n520_), .A3(new_n613_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n549_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n797_), .A2(new_n350_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G169gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT62), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n797_), .A2(new_n848_), .A3(new_n844_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n797_), .B2(new_n844_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n350_), .A2(new_n401_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n847_), .B1(new_n852_), .B2(new_n853_), .ZN(G1348gat));
  INV_X1    g653(.A(new_n852_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n312_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n549_), .B1(new_n781_), .B2(new_n787_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n843_), .A2(new_n368_), .A3(new_n684_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n856_), .A2(new_n368_), .B1(new_n857_), .B2(new_n858_), .ZN(G1349gat));
  NOR3_X1   g658(.A1(new_n852_), .A2(new_n734_), .A3(new_n407_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n640_), .A3(new_n842_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n371_), .B2(new_n861_), .ZN(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n852_), .B2(new_n838_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n619_), .A2(new_n409_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n852_), .B2(new_n864_), .ZN(G1351gat));
  INV_X1    g664(.A(new_n552_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n718_), .A2(new_n564_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n795_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n582_), .B1(new_n869_), .B2(new_n778_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n866_), .B(new_n867_), .C1(new_n870_), .C2(new_n786_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n350_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n312_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g675(.A(new_n734_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT125), .B1(new_n871_), .B2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n828_), .A2(new_n882_), .A3(new_n867_), .A4(new_n877_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT126), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n872_), .A2(new_n882_), .A3(new_n885_), .A4(new_n877_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n881_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n881_), .B1(new_n886_), .B2(new_n884_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1354gat));
  AND3_X1   g688(.A1(new_n872_), .A2(G218gat), .A3(new_n608_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n871_), .A2(new_n602_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n891_), .A2(KEYINPUT127), .ZN(new_n892_));
  AOI21_X1  g691(.A(G218gat), .B1(new_n891_), .B2(KEYINPUT127), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n892_), .B2(new_n893_), .ZN(G1355gat));
endmodule


