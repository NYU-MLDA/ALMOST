//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n994_, new_n995_, new_n997_,
    new_n998_, new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1039_, new_n1040_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1051_, new_n1052_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1065_, new_n1066_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G127gat), .B(G134gat), .Z(new_n204_));
  XOR2_X1   g003(.A(G113gat), .B(G120gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT83), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n204_), .A2(new_n205_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT3), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n217_), .B1(new_n218_), .B2(KEYINPUT1), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT86), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT1), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT87), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n217_), .A2(new_n225_), .A3(KEYINPUT1), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n217_), .B2(KEYINPUT1), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n212_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(G141gat), .B2(G148gat), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n229_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n220_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n211_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n209_), .A2(new_n206_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n220_), .B(new_n238_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n203_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT4), .B1(new_n211_), .B2(new_n236_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n220_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n228_), .A2(new_n233_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT88), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n239_), .B1(new_n246_), .B2(new_n210_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n241_), .B1(new_n247_), .B2(KEYINPUT4), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n240_), .B1(new_n248_), .B2(new_n203_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT0), .ZN(new_n251_));
  INV_X1    g050(.A(G57gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G85gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n259_), .A2(new_n202_), .A3(new_n241_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n260_), .B2(new_n240_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(new_n261_), .A3(KEYINPUT96), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT77), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT77), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(G183gat), .A3(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT78), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT23), .B1(new_n269_), .B2(new_n271_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n268_), .A2(KEYINPUT23), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n268_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n275_), .A2(new_n278_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT25), .B(G183gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(KEYINPUT24), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n288_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(KEYINPUT22), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G169gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n298_), .A3(new_n290_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT22), .B(G169gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT79), .A3(new_n290_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n301_), .A2(new_n303_), .A3(new_n292_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n272_), .B2(KEYINPUT23), .ZN(new_n306_));
  INV_X1    g105(.A(G183gat), .ZN(new_n307_));
  INV_X1    g106(.A(G190gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n285_), .A2(new_n295_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT21), .ZN(new_n312_));
  INV_X1    g111(.A(G204gat), .ZN(new_n313_));
  INV_X1    g112(.A(G197gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT89), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(KEYINPUT89), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G197gat), .A2(G204gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n312_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n312_), .B1(G197gat), .B2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n317_), .A2(new_n318_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n320_), .A2(new_n312_), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n319_), .A2(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT90), .B1(new_n311_), .B2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n282_), .B(new_n281_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n274_), .A2(KEYINPUT78), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n295_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n299_), .A2(new_n300_), .B1(G169gat), .B2(G176gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n310_), .A2(new_n303_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n327_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n328_), .A2(new_n337_), .A3(KEYINPUT20), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n295_), .A2(new_n306_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n283_), .B1(KEYINPUT78), .B2(new_n274_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n343_), .A2(new_n278_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n299_), .A2(new_n292_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n342_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n341_), .B1(new_n346_), .B2(new_n335_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n338_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n328_), .A2(new_n337_), .A3(KEYINPUT20), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT91), .B1(new_n351_), .B2(new_n347_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n285_), .A2(new_n309_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n345_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n354_), .A2(new_n355_), .B1(new_n295_), .B2(new_n306_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(new_n327_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n334_), .B2(new_n335_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n340_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n353_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT97), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n327_), .B1(new_n356_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n346_), .A2(KEYINPUT95), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n340_), .B1(new_n371_), .B2(new_n351_), .ZN(new_n372_));
  OR3_X1    g171(.A1(new_n357_), .A2(new_n340_), .A3(new_n358_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n364_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n367_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT97), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n353_), .A2(new_n377_), .A3(new_n359_), .A4(new_n364_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n366_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n365_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n364_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n367_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n335_), .B1(new_n246_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G228gat), .ZN(new_n387_));
  INV_X1    g186(.A(G233gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n327_), .B1(new_n236_), .B2(KEYINPUT29), .ZN(new_n391_));
  INV_X1    g190(.A(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n390_), .B(new_n393_), .C1(KEYINPUT29), .C2(new_n236_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G22gat), .B(G50gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT28), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n396_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(G15gat), .A2(G43gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G15gat), .A2(G43gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT80), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n407_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n413_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n406_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n331_), .A2(KEYINPUT30), .A3(new_n333_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT30), .B1(new_n331_), .B2(new_n333_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT81), .B(new_n423_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT31), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n288_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n343_), .B2(new_n278_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n301_), .A2(new_n303_), .A3(new_n292_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n432_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n417_), .A2(new_n422_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n331_), .A2(new_n333_), .A3(KEYINPUT30), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT82), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n437_), .A2(new_n438_), .A3(new_n442_), .A4(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n430_), .A2(new_n431_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n431_), .B1(new_n430_), .B2(new_n444_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n211_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n430_), .A2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT31), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n430_), .A2(new_n444_), .A3(new_n431_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n210_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n405_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n211_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n210_), .A3(new_n450_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT84), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n404_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n404_), .A2(new_n454_), .A3(new_n453_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n267_), .B(new_n384_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n455_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n374_), .A2(KEYINPUT32), .A3(new_n364_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n353_), .A2(new_n359_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n262_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n349_), .B1(new_n338_), .B2(new_n348_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n351_), .A2(new_n347_), .A3(KEYINPUT91), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n359_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n375_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n249_), .B2(new_n255_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT33), .B(new_n257_), .C1(new_n260_), .C2(new_n240_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n365_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n247_), .A2(KEYINPUT4), .ZN(new_n472_));
  INV_X1    g271(.A(new_n241_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n255_), .B1(new_n247_), .B2(new_n202_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n474_), .A2(new_n202_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n255_), .B(KEYINPUT93), .C1(new_n247_), .C2(new_n202_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT94), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n476_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n202_), .B1(new_n259_), .B2(new_n241_), .ZN(new_n481_));
  AND4_X1   g280(.A1(KEYINPUT94), .A2(new_n480_), .A3(new_n481_), .A4(new_n478_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n463_), .B1(new_n471_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n459_), .A2(new_n484_), .A3(new_n404_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G1gat), .A2(G8gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT14), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n486_), .A2(new_n487_), .A3(new_n492_), .A4(new_n488_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G43gat), .B(G50gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n499_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510_));
  INV_X1    g309(.A(new_n499_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n497_), .A2(new_n498_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n502_), .A2(KEYINPUT15), .A3(new_n499_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n496_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n516_));
  INV_X1    g315(.A(G141gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G113gat), .ZN(new_n518_));
  INV_X1    g317(.A(G113gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G141gat), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n289_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n520_), .A3(new_n289_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(G197gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n314_), .B1(new_n525_), .B2(new_n521_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n509_), .A2(new_n516_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n509_), .B2(new_n516_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n533_), .B2(KEYINPUT74), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n505_), .A2(new_n507_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n535_), .A2(new_n515_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT75), .B1(new_n534_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n536_), .B2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(KEYINPUT74), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .A4(new_n528_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n458_), .A2(new_n485_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G230gat), .A2(G233gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT64), .Z(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  AND3_X1   g347(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT6), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(KEYINPUT66), .A3(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n557_));
  INV_X1    g356(.A(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n551_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562_));
  INV_X1    g361(.A(G92gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n254_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n562_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n566_), .A2(new_n568_), .A3(KEYINPUT65), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT65), .ZN(new_n570_));
  INV_X1    g369(.A(new_n565_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT9), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n570_), .B1(new_n573_), .B2(new_n567_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n561_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT67), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT65), .B1(new_n566_), .B2(new_n568_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n573_), .A2(new_n570_), .A3(new_n567_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT67), .A3(new_n561_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT68), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n549_), .A2(new_n550_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587_));
  INV_X1    g386(.A(G99gat), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n558_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT68), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n582_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n571_), .A2(new_n572_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT8), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT8), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n551_), .A2(new_n556_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n582_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n596_), .B(new_n593_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n577_), .A2(new_n581_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G71gat), .B(G78gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(G57gat), .B(G64gat), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n601_), .B1(KEYINPUT11), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT11), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n547_), .B1(new_n600_), .B2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n600_), .A2(KEYINPUT12), .A3(new_n606_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n609_));
  INV_X1    g408(.A(new_n593_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n554_), .A2(new_n555_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n598_), .B2(KEYINPUT68), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n612_), .B2(new_n591_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n599_), .B1(new_n613_), .B2(new_n596_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n580_), .A2(KEYINPUT67), .A3(new_n561_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT67), .B1(new_n580_), .B2(new_n561_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n609_), .B1(new_n617_), .B2(new_n605_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n607_), .B1(new_n608_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n605_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n606_), .B(new_n614_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n547_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n625_));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n619_), .A2(new_n623_), .A3(new_n629_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT70), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT70), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n619_), .A2(new_n623_), .A3(new_n633_), .A4(new_n629_), .ZN(new_n634_));
  AOI221_X4 g433(.A(new_n545_), .B1(new_n624_), .B2(new_n630_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n630_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT13), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT71), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT12), .B1(new_n600_), .B2(new_n606_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n617_), .A2(new_n609_), .A3(new_n605_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n642_), .A2(new_n607_), .B1(new_n622_), .B2(new_n547_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n633_), .B1(new_n643_), .B2(new_n629_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n634_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n637_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n545_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT71), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n636_), .A2(KEYINPUT13), .A3(new_n637_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n639_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT36), .Z(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT34), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT35), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n504_), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n617_), .A2(new_n662_), .B1(KEYINPUT35), .B2(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n513_), .A2(new_n514_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n600_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n600_), .A2(new_n504_), .B1(new_n660_), .B2(new_n659_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n661_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n617_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n656_), .B1(new_n666_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n654_), .A2(KEYINPUT36), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n666_), .A2(new_n670_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(KEYINPUT37), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT37), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n666_), .A2(new_n670_), .A3(new_n673_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n671_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(G231gat), .A2(G233gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n496_), .B(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n682_), .A2(new_n606_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(G183gat), .B(G211gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(G127gat), .B(G155gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n686_), .A2(new_n688_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT17), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n682_), .A2(new_n606_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n683_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT17), .ZN(new_n696_));
  INV_X1    g495(.A(new_n691_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n689_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n692_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n683_), .B2(new_n694_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n695_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n651_), .A2(new_n680_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n544_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT98), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n544_), .A2(KEYINPUT98), .A3(new_n703_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n267_), .A2(G1gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT99), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n677_), .A2(new_n671_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n647_), .A2(new_n649_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n534_), .A2(new_n538_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n702_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n379_), .A2(new_n382_), .A3(new_n264_), .A4(new_n265_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n404_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT84), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT84), .B1(new_n453_), .B2(new_n454_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n457_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n459_), .A2(new_n484_), .A3(new_n404_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n714_), .B(new_n717_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n490_), .B1(new_n727_), .B2(new_n266_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT99), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n708_), .A2(new_n730_), .A3(KEYINPUT38), .A4(new_n709_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n712_), .A2(new_n729_), .A3(new_n731_), .ZN(G1324gat));
  NAND4_X1  g531(.A1(new_n706_), .A2(new_n491_), .A3(new_n383_), .A4(new_n707_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n457_), .B1(new_n459_), .B2(new_n719_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n485_), .B1(new_n734_), .B2(new_n718_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n735_), .A2(new_n383_), .A3(new_n714_), .A4(new_n717_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G8gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G8gat), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(KEYINPUT39), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT39), .ZN(new_n741_));
  OAI21_X1  g540(.A(G8gat), .B1(new_n726_), .B2(new_n384_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT100), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n736_), .A2(new_n737_), .A3(G8gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n733_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT40), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT40), .B(new_n733_), .C1(new_n740_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1325gat));
  NOR3_X1   g549(.A1(new_n704_), .A2(G15gat), .A3(new_n459_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT101), .ZN(new_n752_));
  INV_X1    g551(.A(G15gat), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n720_), .A2(new_n721_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n727_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT41), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n756_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n757_), .A3(new_n758_), .ZN(G1326gat));
  OR3_X1    g558(.A1(new_n704_), .A2(G22gat), .A3(new_n404_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G22gat), .B1(new_n726_), .B2(new_n404_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT42), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT42), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(G1327gat));
  NAND2_X1  g563(.A1(new_n539_), .A2(new_n543_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n713_), .A2(new_n702_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n715_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n735_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G29gat), .B1(new_n769_), .B2(new_n266_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n715_), .A2(new_n716_), .A3(new_n701_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n772_));
  XOR2_X1   g571(.A(new_n679_), .B(KEYINPUT103), .Z(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n735_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n680_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n458_), .B2(new_n485_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT44), .B(new_n771_), .C1(new_n774_), .C2(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(G29gat), .A3(new_n266_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n771_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n770_), .B1(new_n779_), .B2(new_n782_), .ZN(G1328gat));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n784_));
  INV_X1    g583(.A(G36gat), .ZN(new_n785_));
  INV_X1    g584(.A(new_n771_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n773_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n772_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n735_), .A2(new_n775_), .A3(new_n680_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n384_), .B1(new_n791_), .B2(KEYINPUT44), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n785_), .B1(new_n792_), .B2(new_n782_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n383_), .A2(new_n785_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT104), .B1(new_n768_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT104), .ZN(new_n796_));
  INV_X1    g595(.A(new_n794_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n544_), .A2(new_n796_), .A3(new_n767_), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n795_), .A2(KEYINPUT45), .A3(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n784_), .B1(new_n793_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n802_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n795_), .B2(new_n798_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n791_), .A2(KEYINPUT44), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n778_), .A2(new_n383_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G36gat), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n810_), .A3(KEYINPUT46), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n804_), .A2(new_n811_), .ZN(G1329gat));
  XNOR2_X1  g611(.A(KEYINPUT105), .B(G43gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n768_), .B2(new_n459_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT106), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT106), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n813_), .C1(new_n768_), .C2(new_n459_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n447_), .A2(new_n451_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n778_), .A2(G43gat), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n820_), .B2(new_n808_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT47), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n818_), .B(new_n823_), .C1(new_n820_), .C2(new_n808_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1330gat));
  AOI21_X1  g624(.A(G50gat), .B1(new_n769_), .B2(new_n719_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n778_), .A2(G50gat), .A3(new_n719_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n782_), .ZN(G1331gat));
  NAND3_X1  g627(.A1(new_n715_), .A2(new_n679_), .A3(new_n701_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT107), .Z(new_n830_));
  INV_X1    g629(.A(new_n716_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n458_), .B2(new_n485_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n252_), .A3(new_n266_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n539_), .A2(new_n701_), .A3(new_n543_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n639_), .A2(new_n650_), .A3(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n837_), .B(new_n714_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT108), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n735_), .A2(KEYINPUT108), .A3(new_n714_), .A4(new_n837_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(new_n266_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n834_), .B1(new_n252_), .B2(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT109), .ZN(G1332gat));
  INV_X1    g643(.A(G64gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n833_), .A2(new_n845_), .A3(new_n383_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n840_), .A2(new_n383_), .A3(new_n841_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT48), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n848_), .A3(G64gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n847_), .B2(G64gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n846_), .B1(new_n849_), .B2(new_n850_), .ZN(G1333gat));
  INV_X1    g650(.A(G71gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n833_), .A2(new_n852_), .A3(new_n754_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n840_), .A2(new_n754_), .A3(new_n841_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(G71gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n854_), .B2(G71gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT110), .B(new_n853_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1334gat));
  INV_X1    g661(.A(G78gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n833_), .A2(new_n863_), .A3(new_n719_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n840_), .A2(new_n719_), .A3(new_n841_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n865_), .A2(new_n866_), .A3(G78gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n865_), .B2(G78gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n867_), .B2(new_n868_), .ZN(G1335gat));
  INV_X1    g668(.A(new_n651_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n766_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(new_n832_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n254_), .A3(new_n266_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n635_), .A2(new_n638_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n831_), .A3(new_n701_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n877_), .A2(new_n266_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n878_), .B2(new_n254_), .ZN(G1336gat));
  NAND3_X1  g678(.A1(new_n872_), .A2(new_n563_), .A3(new_n383_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n877_), .A2(new_n383_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n563_), .ZN(G1337gat));
  NAND2_X1  g681(.A1(new_n877_), .A2(new_n754_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n819_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n883_), .A2(G99gat), .B1(new_n872_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1338gat));
  NAND3_X1  g686(.A1(new_n872_), .A2(new_n558_), .A3(new_n719_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n719_), .B(new_n875_), .C1(new_n774_), .C2(new_n777_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(G106gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n889_), .B2(G106gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n888_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT53), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n895_), .B(new_n888_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1339gat));
  INV_X1    g696(.A(KEYINPUT111), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n835_), .A2(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n539_), .A2(KEYINPUT111), .A3(new_n543_), .A4(new_n701_), .ZN(new_n900_));
  AND4_X1   g699(.A1(new_n675_), .A2(new_n899_), .A3(new_n678_), .A4(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n901_), .A2(new_n647_), .A3(new_n902_), .A4(new_n649_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT112), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n874_), .A2(new_n905_), .A3(new_n902_), .A4(new_n901_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n901_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT54), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n904_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT55), .B(new_n607_), .C1(new_n608_), .C2(new_n618_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n547_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n621_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n914_));
  OAI21_X1  g713(.A(new_n910_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n911_), .B1(new_n642_), .B2(new_n621_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n630_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n630_), .B(new_n918_), .C1(new_n915_), .C2(new_n916_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n716_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n527_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n515_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n528_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n646_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n713_), .B1(new_n923_), .B2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(KEYINPUT57), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT115), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n917_), .A2(KEYINPUT56), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n934_), .B(new_n630_), .C1(new_n915_), .C2(new_n916_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n927_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(KEYINPUT58), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n679_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n939_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n933_), .A2(new_n941_), .A3(new_n936_), .A4(new_n935_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(KEYINPUT57), .A2(new_n930_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT115), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(new_n930_), .B2(KEYINPUT57), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n932_), .A2(new_n943_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n909_), .B1(new_n946_), .B2(new_n702_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n384_), .A2(new_n266_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n723_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n947_), .A2(new_n950_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n951_), .A2(new_n519_), .A3(new_n831_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n923_), .A2(new_n929_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n953_), .A2(KEYINPUT57), .A3(new_n714_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n935_), .A2(new_n636_), .A3(new_n928_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n642_), .A2(new_n621_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n547_), .ZN(new_n957_));
  OAI211_X1 g756(.A(new_n957_), .B(new_n910_), .C1(new_n913_), .C2(new_n914_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n934_), .B1(new_n958_), .B2(new_n630_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n939_), .B1(new_n955_), .B2(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n960_), .A2(new_n680_), .A3(new_n942_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n954_), .A2(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n702_), .B1(new_n962_), .B2(new_n931_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n909_), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  OAI211_X1 g764(.A(KEYINPUT118), .B(new_n702_), .C1(new_n962_), .C2(new_n931_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  XOR2_X1   g766(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n968_));
  NAND3_X1  g767(.A1(new_n967_), .A2(new_n949_), .A3(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(KEYINPUT59), .B1(new_n947_), .B2(new_n950_), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n969_), .A2(new_n765_), .A3(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n952_), .B1(new_n971_), .B2(new_n519_), .ZN(G1340gat));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n973_), .B1(new_n874_), .B2(G120gat), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n946_), .A2(new_n702_), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n949_), .B(new_n974_), .C1(new_n975_), .C2(new_n909_), .ZN(new_n976_));
  NAND4_X1  g775(.A1(new_n969_), .A2(new_n976_), .A3(new_n651_), .A4(new_n970_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n977_), .A2(G120gat), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n978_), .B1(KEYINPUT60), .B2(new_n976_), .ZN(G1341gat));
  INV_X1    g778(.A(G127gat), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n951_), .A2(new_n980_), .A3(new_n701_), .ZN(new_n981_));
  AND3_X1   g780(.A1(new_n969_), .A2(new_n701_), .A3(new_n970_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n982_), .B2(new_n980_), .ZN(G1342gat));
  INV_X1    g782(.A(G134gat), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n951_), .A2(new_n984_), .A3(new_n713_), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n969_), .A2(new_n680_), .A3(new_n970_), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n985_), .B1(new_n986_), .B2(new_n984_), .ZN(G1343gat));
  NOR2_X1   g786(.A1(new_n948_), .A2(new_n722_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(KEYINPUT119), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n947_), .A2(new_n989_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n990_), .A2(new_n831_), .ZN(new_n991_));
  XNOR2_X1  g790(.A(KEYINPUT120), .B(G141gat), .ZN(new_n992_));
  XOR2_X1   g791(.A(new_n991_), .B(new_n992_), .Z(G1344gat));
  NAND2_X1  g792(.A1(new_n990_), .A2(new_n651_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(KEYINPUT121), .B(G148gat), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n994_), .B(new_n995_), .ZN(G1345gat));
  NAND2_X1  g795(.A1(new_n990_), .A2(new_n701_), .ZN(new_n997_));
  XNOR2_X1  g796(.A(KEYINPUT61), .B(G155gat), .ZN(new_n998_));
  XNOR2_X1  g797(.A(new_n997_), .B(new_n998_), .ZN(G1346gat));
  AOI21_X1  g798(.A(G162gat), .B1(new_n990_), .B2(new_n713_), .ZN(new_n1000_));
  AND2_X1   g799(.A1(new_n773_), .A2(G162gat), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n1000_), .B1(new_n990_), .B2(new_n1001_), .ZN(G1347gat));
  NAND3_X1  g801(.A1(new_n754_), .A2(new_n267_), .A3(new_n383_), .ZN(new_n1003_));
  AND2_X1   g802(.A1(new_n1003_), .A2(KEYINPUT122), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(new_n1003_), .A2(KEYINPUT122), .ZN(new_n1005_));
  OAI21_X1  g804(.A(new_n404_), .B1(new_n1004_), .B2(new_n1005_), .ZN(new_n1006_));
  AOI211_X1 g805(.A(new_n716_), .B(new_n1006_), .C1(new_n965_), .C2(new_n966_), .ZN(new_n1007_));
  OAI21_X1  g806(.A(KEYINPUT123), .B1(new_n1007_), .B2(new_n289_), .ZN(new_n1008_));
  INV_X1    g807(.A(new_n1006_), .ZN(new_n1009_));
  NAND3_X1  g808(.A1(new_n904_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n1010_));
  OR2_X1    g809(.A1(new_n930_), .A2(KEYINPUT57), .ZN(new_n1011_));
  AOI21_X1  g810(.A(new_n701_), .B1(new_n943_), .B2(new_n1011_), .ZN(new_n1012_));
  OAI21_X1  g811(.A(new_n1010_), .B1(new_n1012_), .B2(KEYINPUT118), .ZN(new_n1013_));
  INV_X1    g812(.A(new_n966_), .ZN(new_n1014_));
  OAI211_X1 g813(.A(new_n831_), .B(new_n1009_), .C1(new_n1013_), .C2(new_n1014_), .ZN(new_n1015_));
  INV_X1    g814(.A(KEYINPUT123), .ZN(new_n1016_));
  NAND3_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .A3(G169gat), .ZN(new_n1017_));
  NAND3_X1  g816(.A1(new_n1008_), .A2(KEYINPUT62), .A3(new_n1017_), .ZN(new_n1018_));
  AND4_X1   g817(.A1(new_n831_), .A2(new_n967_), .A3(new_n302_), .A4(new_n1009_), .ZN(new_n1019_));
  AOI21_X1  g818(.A(new_n1016_), .B1(new_n1015_), .B2(G169gat), .ZN(new_n1020_));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1021_));
  AOI21_X1  g820(.A(new_n1019_), .B1(new_n1020_), .B2(new_n1021_), .ZN(new_n1022_));
  NAND2_X1  g821(.A1(new_n1018_), .A2(new_n1022_), .ZN(G1348gat));
  NAND2_X1  g822(.A1(new_n967_), .A2(new_n1009_), .ZN(new_n1024_));
  INV_X1    g823(.A(new_n1024_), .ZN(new_n1025_));
  AOI21_X1  g824(.A(G176gat), .B1(new_n1025_), .B2(new_n715_), .ZN(new_n1026_));
  NOR2_X1   g825(.A1(new_n947_), .A2(new_n719_), .ZN(new_n1027_));
  NOR2_X1   g826(.A1(new_n1004_), .A2(new_n1005_), .ZN(new_n1028_));
  NOR3_X1   g827(.A1(new_n1028_), .A2(new_n290_), .A3(new_n870_), .ZN(new_n1029_));
  AOI21_X1  g828(.A(new_n1026_), .B1(new_n1027_), .B2(new_n1029_), .ZN(G1349gat));
  OAI211_X1 g829(.A(new_n1027_), .B(new_n701_), .C1(new_n1005_), .C2(new_n1004_), .ZN(new_n1031_));
  NAND2_X1  g830(.A1(new_n1031_), .A2(new_n307_), .ZN(new_n1032_));
  NOR2_X1   g831(.A1(new_n702_), .A2(new_n286_), .ZN(new_n1033_));
  NAND3_X1  g832(.A1(new_n1025_), .A2(KEYINPUT124), .A3(new_n1033_), .ZN(new_n1034_));
  INV_X1    g833(.A(KEYINPUT124), .ZN(new_n1035_));
  INV_X1    g834(.A(new_n1033_), .ZN(new_n1036_));
  OAI21_X1  g835(.A(new_n1035_), .B1(new_n1024_), .B2(new_n1036_), .ZN(new_n1037_));
  AND3_X1   g836(.A1(new_n1032_), .A2(new_n1034_), .A3(new_n1037_), .ZN(G1350gat));
  OAI21_X1  g837(.A(G190gat), .B1(new_n1024_), .B2(new_n679_), .ZN(new_n1039_));
  NAND2_X1  g838(.A1(new_n713_), .A2(new_n287_), .ZN(new_n1040_));
  OAI21_X1  g839(.A(new_n1039_), .B1(new_n1024_), .B2(new_n1040_), .ZN(G1351gat));
  NOR3_X1   g840(.A1(new_n722_), .A2(new_n384_), .A3(new_n266_), .ZN(new_n1042_));
  OAI21_X1  g841(.A(new_n1042_), .B1(new_n975_), .B2(new_n909_), .ZN(new_n1043_));
  OAI211_X1 g842(.A(KEYINPUT125), .B(new_n314_), .C1(new_n1043_), .C2(new_n716_), .ZN(new_n1044_));
  INV_X1    g843(.A(KEYINPUT125), .ZN(new_n1045_));
  INV_X1    g844(.A(new_n1042_), .ZN(new_n1046_));
  NOR3_X1   g845(.A1(new_n947_), .A2(new_n716_), .A3(new_n1046_), .ZN(new_n1047_));
  OAI21_X1  g846(.A(new_n1045_), .B1(new_n1047_), .B2(G197gat), .ZN(new_n1048_));
  NAND2_X1  g847(.A1(new_n1047_), .A2(G197gat), .ZN(new_n1049_));
  AND3_X1   g848(.A1(new_n1044_), .A2(new_n1048_), .A3(new_n1049_), .ZN(G1352gat));
  NOR2_X1   g849(.A1(new_n947_), .A2(new_n1046_), .ZN(new_n1051_));
  NAND2_X1  g850(.A1(new_n1051_), .A2(new_n651_), .ZN(new_n1052_));
  XNOR2_X1  g851(.A(new_n1052_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g852(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1054_));
  INV_X1    g853(.A(KEYINPUT63), .ZN(new_n1055_));
  INV_X1    g854(.A(G211gat), .ZN(new_n1056_));
  NOR2_X1   g855(.A1(new_n1055_), .A2(new_n1056_), .ZN(new_n1057_));
  NOR4_X1   g856(.A1(new_n1043_), .A2(new_n702_), .A3(new_n1054_), .A4(new_n1057_), .ZN(new_n1058_));
  INV_X1    g857(.A(KEYINPUT126), .ZN(new_n1059_));
  NOR2_X1   g858(.A1(new_n1043_), .A2(new_n702_), .ZN(new_n1060_));
  NAND2_X1  g859(.A1(new_n1055_), .A2(new_n1056_), .ZN(new_n1061_));
  OAI21_X1  g860(.A(new_n1059_), .B1(new_n1060_), .B2(new_n1061_), .ZN(new_n1062_));
  OAI211_X1 g861(.A(KEYINPUT126), .B(new_n1054_), .C1(new_n1043_), .C2(new_n702_), .ZN(new_n1063_));
  AOI21_X1  g862(.A(new_n1058_), .B1(new_n1062_), .B2(new_n1063_), .ZN(G1354gat));
  OR3_X1    g863(.A1(new_n1043_), .A2(G218gat), .A3(new_n714_), .ZN(new_n1065_));
  OAI21_X1  g864(.A(G218gat), .B1(new_n1043_), .B2(new_n679_), .ZN(new_n1066_));
  NAND2_X1  g865(.A1(new_n1065_), .A2(new_n1066_), .ZN(G1355gat));
endmodule


