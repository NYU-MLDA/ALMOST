//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n987_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT22), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT81), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n221_), .B2(KEYINPUT23), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n215_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT26), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G190gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT23), .B1(new_n218_), .B2(new_n220_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT78), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(G169gat), .B2(G176gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT24), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  NOR3_X1   g041(.A1(new_n233_), .A2(new_n237_), .A3(new_n242_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n239_), .A2(new_n241_), .A3(KEYINPUT24), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(KEYINPUT80), .A3(new_n207_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n241_), .A3(KEYINPUT24), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n206_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n223_), .B1(new_n243_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT82), .B(G15gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n250_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G127gat), .B(G134gat), .Z(new_n255_));
  INV_X1    g054(.A(G120gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G113gat), .ZN(new_n257_));
  INV_X1    g056(.A(G113gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G120gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n254_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G71gat), .B(G99gat), .ZN(new_n267_));
  INV_X1    g066(.A(G43gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT30), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n266_), .A2(new_n271_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT83), .B1(new_n277_), .B2(KEYINPUT1), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(G155gat), .A4(G162gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(KEYINPUT1), .ZN(new_n282_));
  OR2_X1    g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G141gat), .B(G148gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n277_), .A3(new_n283_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n264_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n276_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT91), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n264_), .A2(new_n296_), .A3(new_n286_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(new_n297_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n302_), .B2(KEYINPUT4), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n286_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n265_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n264_), .A2(new_n296_), .A3(new_n286_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n305_), .A2(new_n300_), .A3(KEYINPUT4), .A4(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n299_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n306_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n276_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT92), .B(G85gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT0), .B(G57gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n299_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT91), .B1(new_n310_), .B2(new_n298_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(new_n307_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n323_), .B2(new_n312_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n275_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT99), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT18), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G204gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT85), .B1(new_n338_), .B2(G197gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n340_));
  INV_X1    g139(.A(G197gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(G204gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(G197gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n339_), .A2(new_n342_), .A3(new_n336_), .A4(new_n343_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(new_n335_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT84), .B1(new_n348_), .B2(new_n336_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(G204gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n343_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT21), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n347_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n347_), .B2(new_n354_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n345_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n215_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n204_), .A2(new_n360_), .A3(new_n205_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n206_), .A2(KEYINPUT89), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n359_), .A2(new_n213_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n244_), .A2(new_n202_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n226_), .A2(new_n231_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n365_), .A2(new_n224_), .B1(new_n366_), .B2(new_n238_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n222_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n358_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n345_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n352_), .B1(new_n351_), .B2(KEYINPUT21), .ZN(new_n372_));
  AOI211_X1 g171(.A(KEYINPUT84), .B(new_n336_), .C1(new_n350_), .C2(new_n343_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n346_), .A2(new_n335_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT86), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n347_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n371_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n250_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT19), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n370_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n358_), .B2(new_n369_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n376_), .A2(new_n377_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n250_), .A2(new_n386_), .A3(new_n345_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n383_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n334_), .B1(new_n382_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n369_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT20), .B1(new_n378_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n222_), .A2(new_n215_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(new_n207_), .A3(new_n213_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n245_), .A2(new_n248_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n239_), .A2(new_n241_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n366_), .ZN(new_n396_));
  OAI221_X1 g195(.A(new_n396_), .B1(new_n234_), .B2(new_n236_), .C1(new_n232_), .C2(new_n229_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n358_), .A2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n381_), .B1(new_n391_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n384_), .B1(new_n378_), .B2(new_n390_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n358_), .A2(new_n398_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n383_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n333_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n389_), .A2(KEYINPUT90), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT90), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n400_), .A2(new_n403_), .A3(new_n407_), .A4(new_n333_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n381_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT95), .B(new_n381_), .C1(new_n370_), .C2(new_n379_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n358_), .A2(new_n369_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n387_), .A3(KEYINPUT20), .A4(new_n383_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT96), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n385_), .A2(new_n418_), .A3(new_n383_), .A4(new_n387_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n413_), .A2(new_n414_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n410_), .B1(new_n420_), .B2(new_n333_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n409_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT98), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n409_), .A2(new_n421_), .A3(KEYINPUT98), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427_));
  INV_X1    g226(.A(G228gat), .ZN(new_n428_));
  INV_X1    g227(.A(G233gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n304_), .A2(KEYINPUT29), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n358_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n358_), .B2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n427_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G22gat), .B(G50gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n304_), .A2(KEYINPUT29), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n444_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n442_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n442_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n449_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n437_), .A2(KEYINPUT87), .A3(new_n433_), .A4(new_n438_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n441_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT88), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n436_), .A2(new_n452_), .A3(new_n439_), .A4(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n329_), .B1(new_n426_), .B2(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n409_), .A2(new_n421_), .A3(KEYINPUT98), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT98), .B1(new_n409_), .B2(new_n421_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n329_), .B(new_n461_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n328_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT97), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n309_), .A2(KEYINPUT33), .A3(new_n313_), .A4(new_n318_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT93), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n319_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n322_), .A2(new_n307_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n312_), .B1(new_n473_), .B2(new_n299_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT33), .A4(new_n318_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n473_), .B(new_n276_), .C1(KEYINPUT4), .C2(new_n305_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n320_), .B1(new_n310_), .B2(new_n276_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n470_), .A2(new_n472_), .A3(new_n476_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n405_), .A2(new_n408_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n420_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n400_), .A2(new_n487_), .A3(new_n403_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n325_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n484_), .A2(new_n485_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n468_), .B1(new_n493_), .B2(new_n460_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n483_), .B1(new_n408_), .B2(new_n405_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT97), .B(new_n461_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n460_), .A2(new_n326_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n422_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n275_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n467_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT74), .B(G8gat), .ZN(new_n512_));
  INV_X1    g311(.A(G1gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n511_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n511_), .B(new_n517_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n510_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n510_), .A3(new_n520_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT76), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n525_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n506_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n509_), .B(KEYINPUT15), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n520_), .A3(new_n519_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(new_n522_), .A3(new_n505_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G169gat), .B(G197gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n522_), .A2(KEYINPUT76), .A3(new_n523_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n526_), .B1(new_n525_), .B2(new_n521_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n505_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n531_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n536_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n519_), .A2(new_n520_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT75), .ZN(new_n544_));
  AND2_X1   g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(KEYINPUT11), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551_));
  INV_X1    g350(.A(G64gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(G57gat), .ZN(new_n553_));
  INV_X1    g352(.A(G57gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G64gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n555_), .A3(KEYINPUT11), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n550_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n547_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n547_), .A2(new_n559_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT16), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n560_), .A2(new_n561_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n559_), .A2(KEYINPUT66), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT66), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n570_), .B(new_n550_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n547_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n569_), .A2(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n546_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n565_), .B(KEYINPUT17), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n568_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT36), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT6), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592_));
  INV_X1    g391(.A(G99gat), .ZN(new_n593_));
  INV_X1    g392(.A(G106gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n588_), .B1(new_n591_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT8), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT8), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n600_), .B(new_n588_), .C1(new_n591_), .C2(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT64), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(KEYINPUT64), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n594_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n591_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n587_), .B1(new_n586_), .B2(KEYINPUT9), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n585_), .A2(KEYINPUT65), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT65), .B1(new_n585_), .B2(new_n613_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n602_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n618_), .A2(new_n529_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n591_), .B1(new_n609_), .B2(new_n594_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n616_), .A2(new_n624_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(KEYINPUT72), .A3(new_n509_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT72), .B1(new_n625_), .B2(new_n509_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n622_), .A2(new_n619_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI221_X1 g429(.A(new_n623_), .B1(new_n619_), .B2(new_n622_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n584_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT73), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n630_), .A2(new_n631_), .A3(KEYINPUT73), .A4(new_n633_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n579_), .B(new_n632_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n637_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n632_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n579_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n578_), .A2(new_n639_), .A3(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT5), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n646_), .B(new_n647_), .Z(new_n648_));
  NAND4_X1  g447(.A1(new_n602_), .A2(new_n617_), .A3(new_n571_), .A4(new_n569_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT67), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT67), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n574_), .A2(new_n625_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n618_), .A2(new_n572_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT68), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT12), .B1(new_n618_), .B2(new_n572_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT12), .B(new_n550_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n618_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n660_), .A2(new_n656_), .A3(new_n649_), .A4(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n655_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n648_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n654_), .A2(new_n657_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT68), .ZN(new_n669_));
  INV_X1    g468(.A(new_n648_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n664_), .A3(new_n658_), .A4(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n667_), .A2(KEYINPUT69), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT69), .B1(new_n667_), .B2(new_n671_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n674_));
  OR3_X1    g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n644_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n504_), .A2(new_n542_), .A3(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n679_), .A2(G1gat), .A3(new_n326_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n680_), .A2(KEYINPUT38), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n677_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n542_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n568_), .A2(new_n577_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT99), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n327_), .B1(new_n688_), .B2(new_n465_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n461_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n499_), .B1(new_n690_), .B2(new_n468_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n275_), .B1(new_n691_), .B2(new_n497_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n686_), .B(new_n642_), .C1(new_n689_), .C2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G1gat), .B1(new_n693_), .B2(new_n326_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n681_), .A2(new_n682_), .A3(new_n694_), .ZN(G1324gat));
  OAI21_X1  g494(.A(G8gat), .B1(new_n693_), .B2(new_n426_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT39), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT39), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(G8gat), .C1(new_n693_), .C2(new_n426_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n679_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n426_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n512_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT101), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n700_), .A2(new_n706_), .A3(new_n703_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n705_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1325gat));
  OAI21_X1  g510(.A(G15gat), .B1(new_n693_), .B2(new_n502_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT41), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n679_), .A2(G15gat), .A3(new_n502_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1326gat));
  OAI21_X1  g514(.A(G22gat), .B1(new_n693_), .B2(new_n461_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n461_), .A2(G22gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n679_), .B2(new_n719_), .ZN(G1327gat));
  AOI21_X1  g519(.A(new_n632_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n685_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT104), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n683_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n504_), .A2(new_n542_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n726_), .B2(new_n325_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n639_), .A2(new_n643_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n728_), .B(new_n729_), .C1(new_n689_), .C2(new_n692_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n728_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n467_), .B2(new_n503_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n729_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n684_), .A2(new_n578_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(KEYINPUT44), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n736_), .B2(new_n737_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n325_), .A2(G29gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n727_), .B1(new_n740_), .B2(new_n741_), .ZN(G1328gat));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n743_), .A3(new_n702_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT45), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n738_), .A2(new_n739_), .A3(new_n426_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n743_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n745_), .B(new_n748_), .C1(new_n743_), .C2(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1329gat));
  NOR2_X1   g551(.A1(new_n502_), .A2(new_n268_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n740_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n268_), .B1(new_n725_), .B2(new_n502_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT106), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1330gat));
  NOR3_X1   g561(.A1(new_n738_), .A2(new_n739_), .A3(new_n461_), .ZN(new_n763_));
  INV_X1    g562(.A(G50gat), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n460_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT108), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n763_), .A2(new_n764_), .B1(new_n725_), .B2(new_n766_), .ZN(G1331gat));
  AOI21_X1  g566(.A(new_n721_), .B1(new_n467_), .B2(new_n503_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n683_), .A2(new_n542_), .A3(new_n685_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n770_), .A2(new_n554_), .A3(new_n326_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772_));
  INV_X1    g571(.A(new_n542_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n504_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n504_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n683_), .A2(new_n644_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT109), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n554_), .B1(new_n781_), .B2(new_n326_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n782_), .A2(KEYINPUT111), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(KEYINPUT111), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n771_), .B1(new_n783_), .B2(new_n784_), .ZN(G1332gat));
  INV_X1    g584(.A(new_n770_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n552_), .B1(new_n786_), .B2(new_n702_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n787_), .A2(new_n788_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n702_), .A2(new_n552_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n790_), .A2(new_n791_), .B1(new_n781_), .B2(new_n792_), .ZN(G1333gat));
  OAI21_X1  g592(.A(G71gat), .B1(new_n770_), .B2(new_n502_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT49), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n502_), .A2(G71gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n781_), .B2(new_n796_), .ZN(G1334gat));
  OAI21_X1  g596(.A(G78gat), .B1(new_n770_), .B2(new_n461_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT50), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n461_), .A2(G78gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n781_), .B2(new_n800_), .ZN(G1335gat));
  INV_X1    g600(.A(new_n683_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n723_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n325_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n683_), .A2(new_n542_), .A3(new_n578_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n736_), .A2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT112), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n325_), .A2(G85gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(G1336gat));
  AOI21_X1  g609(.A(G92gat), .B1(new_n804_), .B2(new_n702_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n702_), .A2(G92gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n808_), .B2(new_n812_), .ZN(G1337gat));
  NAND3_X1  g612(.A1(new_n804_), .A2(new_n275_), .A3(new_n609_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G99gat), .B1(new_n807_), .B2(new_n502_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n736_), .A2(new_n460_), .A3(new_n806_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(G106gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n818_), .B2(G106gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n806_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n728_), .B1(new_n689_), .B2(new_n692_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n735_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n461_), .B(new_n824_), .C1(new_n827_), .C2(new_n730_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT114), .B(new_n822_), .C1(new_n828_), .C2(new_n594_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n804_), .A2(new_n594_), .A3(new_n460_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT53), .B1(new_n823_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT114), .B1(new_n828_), .B2(new_n594_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n818_), .A2(new_n819_), .A3(G106gat), .ZN(new_n834_));
  INV_X1    g633(.A(new_n822_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n829_), .A4(new_n830_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n838_), .ZN(G1339gat));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n678_), .A2(KEYINPUT115), .A3(new_n840_), .A4(new_n773_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n721_), .A2(KEYINPUT37), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n842_), .A2(new_n685_), .A3(new_n638_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n683_), .A2(new_n840_), .A3(new_n773_), .A4(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n683_), .A2(new_n773_), .A3(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n841_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n671_), .A2(new_n542_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n671_), .A2(KEYINPUT116), .A3(new_n542_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n663_), .A2(new_n649_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n657_), .B1(new_n856_), .B2(new_n659_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT55), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n664_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n856_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n857_), .A3(KEYINPUT55), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT56), .B1(new_n862_), .B2(new_n648_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n864_), .B(new_n670_), .C1(new_n859_), .C2(new_n861_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n854_), .B(new_n855_), .C1(new_n863_), .C2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n861_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n860_), .B1(KEYINPUT55), .B2(new_n857_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n648_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n864_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n862_), .A2(KEYINPUT56), .A3(new_n648_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n874_), .A2(KEYINPUT117), .A3(new_n854_), .A4(new_n855_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n672_), .A2(new_n673_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n505_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n521_), .A2(new_n505_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n534_), .B1(new_n530_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n535_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n868_), .A2(new_n875_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n851_), .B1(new_n883_), .B2(new_n642_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n874_), .A2(new_n881_), .A3(new_n671_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n874_), .A2(new_n881_), .A3(KEYINPUT58), .A4(new_n671_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n728_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n884_), .B2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n883_), .A2(KEYINPUT57), .A3(new_n642_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n866_), .A2(new_n867_), .B1(new_n876_), .B2(new_n881_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n721_), .B1(new_n894_), .B2(new_n875_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n893_), .B(new_n889_), .C1(new_n895_), .C2(new_n851_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n891_), .A2(new_n892_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n849_), .B1(new_n897_), .B2(new_n685_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n688_), .A2(new_n465_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n502_), .A2(new_n326_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n901_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n892_), .B(new_n889_), .C1(new_n895_), .C2(new_n851_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n685_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n841_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  OAI22_X1  g706(.A1(new_n898_), .A2(new_n902_), .B1(new_n907_), .B2(new_n900_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G113gat), .B1(new_n908_), .B2(new_n773_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n258_), .A3(new_n542_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1340gat));
  OAI21_X1  g710(.A(G120gat), .B1(new_n908_), .B2(new_n683_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n907_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n256_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(KEYINPUT60), .B2(new_n256_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n912_), .B1(new_n913_), .B2(new_n915_), .ZN(G1341gat));
  OAI21_X1  g715(.A(G127gat), .B1(new_n908_), .B2(new_n685_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n685_), .A2(G127gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n913_), .B2(new_n918_), .ZN(G1342gat));
  OAI21_X1  g718(.A(G134gat), .B1(new_n908_), .B2(new_n731_), .ZN(new_n920_));
  OR3_X1    g719(.A1(new_n913_), .A2(G134gat), .A3(new_n642_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT120), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n920_), .A2(new_n924_), .A3(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1343gat));
  NAND4_X1  g725(.A1(new_n426_), .A2(new_n502_), .A3(new_n460_), .A4(new_n325_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT121), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n542_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n802_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n578_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1346gat));
  AOI21_X1  g735(.A(G162gat), .B1(new_n929_), .B2(new_n721_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n728_), .A2(G162gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT122), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n929_), .B2(new_n939_), .ZN(G1347gat));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n426_), .A2(new_n460_), .A3(new_n327_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n898_), .A2(new_n773_), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945_));
  OAI21_X1  g744(.A(G169gat), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n897_), .A2(new_n685_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n542_), .B(new_n942_), .C1(new_n947_), .C2(new_n849_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(KEYINPUT123), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n941_), .B1(new_n946_), .B2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n208_), .B1(new_n948_), .B2(KEYINPUT123), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n944_), .A2(new_n945_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n951_), .A2(KEYINPUT62), .A3(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n944_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n950_), .A2(new_n953_), .A3(new_n954_), .ZN(G1348gat));
  AOI21_X1  g754(.A(new_n943_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n956_), .A2(G176gat), .A3(new_n802_), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT124), .Z(new_n958_));
  NOR2_X1   g757(.A1(new_n898_), .A2(new_n943_), .ZN(new_n959_));
  AOI21_X1  g758(.A(G176gat), .B1(new_n959_), .B2(new_n802_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n958_), .A2(new_n960_), .ZN(G1349gat));
  NOR2_X1   g760(.A1(new_n685_), .A2(new_n224_), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n959_), .A2(KEYINPUT125), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n959_), .B2(new_n962_), .ZN(new_n964_));
  AOI21_X1  g763(.A(G183gat), .B1(new_n956_), .B2(new_n578_), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n959_), .A2(new_n365_), .A3(new_n721_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n898_), .A2(new_n731_), .A3(new_n943_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n968_), .B2(new_n225_), .ZN(G1351gat));
  NAND2_X1  g768(.A1(new_n905_), .A2(new_n906_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n426_), .A2(new_n275_), .A3(new_n498_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n972_), .A2(new_n773_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT126), .B(G197gat), .Z(new_n974_));
  XNOR2_X1  g773(.A(new_n973_), .B(new_n974_), .ZN(G1352gat));
  NOR2_X1   g774(.A1(new_n972_), .A2(new_n683_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(new_n338_), .ZN(G1353gat));
  INV_X1    g776(.A(new_n972_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(new_n578_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  AND2_X1   g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  NOR3_X1   g780(.A1(new_n979_), .A2(new_n980_), .A3(new_n981_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n982_), .B1(new_n979_), .B2(new_n980_), .ZN(G1354gat));
  AND3_X1   g782(.A1(new_n978_), .A2(G218gat), .A3(new_n728_), .ZN(new_n984_));
  NOR3_X1   g783(.A1(new_n972_), .A2(KEYINPUT127), .A3(new_n642_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n985_), .A2(G218gat), .ZN(new_n986_));
  OAI21_X1  g785(.A(KEYINPUT127), .B1(new_n972_), .B2(new_n642_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n984_), .B1(new_n986_), .B2(new_n987_), .ZN(G1355gat));
endmodule


