//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G85gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT6), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n209_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT8), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n208_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n214_), .B1(new_n219_), .B2(new_n205_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n210_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n215_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n205_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n214_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n212_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT66), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(new_n212_), .C1(new_n220_), .C2(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT12), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n231_), .A2(new_n232_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n239_), .B(KEYINPUT69), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n227_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT12), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n228_), .A2(new_n239_), .A3(new_n230_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n245_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G120gat), .B(G148gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT5), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G176gat), .B(G204gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n248_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n228_), .A2(new_n257_), .A3(new_n239_), .A4(new_n230_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n228_), .A2(new_n230_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n239_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n246_), .A2(KEYINPUT67), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n256_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n246_), .A2(KEYINPUT67), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n265_), .B(new_n258_), .C1(new_n239_), .C2(new_n259_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n266_), .B2(new_n256_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n251_), .B(new_n255_), .C1(new_n264_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT13), .ZN(new_n269_));
  INV_X1    g068(.A(new_n251_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n262_), .A2(new_n263_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(KEYINPUT68), .A3(new_n256_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n255_), .B(KEYINPUT71), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n268_), .B(new_n269_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n251_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n269_), .B1(new_n279_), .B2(new_n268_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G29gat), .B(G36gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G43gat), .B(G50gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n288_), .B(new_n291_), .Z(new_n292_));
  NAND2_X1  g091(.A1(G229gat), .A2(G233gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n291_), .B(KEYINPUT15), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n288_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n288_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n297_), .B2(new_n291_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n292_), .A2(new_n294_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G141gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G169gat), .B(G197gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n300_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT79), .B1(new_n299_), .B2(new_n304_), .ZN(new_n307_));
  OAI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n297_), .B(new_n239_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G127gat), .B(G155gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G183gat), .B(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT17), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n312_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n312_), .A2(new_n320_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n281_), .A2(new_n309_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(G197gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336_));
  INV_X1    g135(.A(G197gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(G204gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n345_));
  INV_X1    g144(.A(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n337_), .A2(G204gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n334_), .A2(G197gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n337_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n346_), .B1(new_n352_), .B2(KEYINPUT21), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n338_), .A2(new_n339_), .ZN(new_n355_));
  AND4_X1   g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n341_), .A4(new_n347_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n345_), .B(new_n353_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n334_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT87), .B1(new_n334_), .B2(G197gat), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n341_), .B(new_n347_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT88), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n340_), .A2(new_n354_), .A3(new_n341_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n345_), .B1(new_n365_), .B2(new_n353_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n344_), .B1(new_n359_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n368_), .A2(KEYINPUT90), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(KEYINPUT90), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n376_));
  INV_X1    g175(.A(G169gat), .ZN(new_n377_));
  INV_X1    g176(.A(G176gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n379_), .A2(KEYINPUT24), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT23), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n387_));
  AND4_X1   g186(.A1(new_n375_), .A2(new_n382_), .A3(new_n385_), .A4(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n374_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n373_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n389_), .B1(new_n374_), .B2(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n381_), .A2(KEYINPUT91), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n381_), .A2(KEYINPUT91), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT22), .B(G169gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n378_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n372_), .A2(new_n388_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n333_), .B1(new_n367_), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT89), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n343_), .B1(new_n402_), .B2(new_n358_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT82), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G169gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n404_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n377_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n385_), .A2(new_n392_), .A3(new_n375_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n379_), .A2(new_n380_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n386_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n370_), .A2(new_n368_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n391_), .A2(new_n413_), .A3(new_n382_), .A4(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n403_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n332_), .B1(new_n400_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n332_), .B1(new_n403_), .B2(new_n417_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n344_), .B(new_n398_), .C1(new_n359_), .C2(new_n366_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT20), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n329_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT0), .B(G57gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G113gat), .B(G120gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT84), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436_));
  INV_X1    g235(.A(G141gat), .ZN(new_n437_));
  INV_X1    g236(.A(G148gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G141gat), .A2(G148gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT2), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n435_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n437_), .A2(new_n438_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n440_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT1), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n446_), .B(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n435_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n433_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n435_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n432_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT92), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n429_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n456_), .A3(KEYINPUT4), .ZN(new_n461_));
  INV_X1    g260(.A(new_n458_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n433_), .B(new_n463_), .C1(new_n447_), .C2(new_n452_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT33), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n458_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n428_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT20), .B1(new_n403_), .B2(new_n398_), .ZN(new_n472_));
  AOI211_X1 g271(.A(new_n343_), .B(new_n416_), .C1(new_n402_), .C2(new_n358_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n331_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n329_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n331_), .B1(new_n367_), .B2(new_n416_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n333_), .B1(new_n403_), .B2(new_n398_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT33), .B(new_n428_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n424_), .A2(new_n471_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n461_), .A2(new_n464_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n458_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n469_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n429_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n470_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n475_), .A2(KEYINPUT32), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n488_), .A2(new_n474_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n488_), .B2(new_n474_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n486_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n367_), .A2(new_n416_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(new_n477_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n422_), .A2(KEYINPUT94), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n331_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n472_), .A2(new_n331_), .A3(new_n473_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n493_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n481_), .B1(new_n492_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n447_), .A2(new_n452_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n403_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n507_), .A2(new_n511_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n505_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT28), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(KEYINPUT28), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G22gat), .B(G50gat), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n515_), .A2(KEYINPUT28), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(new_n516_), .ZN(new_n523_));
  OAI22_X1  g322(.A1(new_n513_), .A2(new_n514_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n520_), .A2(new_n523_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n403_), .A2(new_n506_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n510_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n527_), .A3(new_n512_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n502_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT96), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n419_), .A2(new_n423_), .A3(new_n329_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n475_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n486_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n479_), .A2(KEYINPUT27), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n498_), .A2(new_n500_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n540_), .B2(new_n329_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n532_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n477_), .A2(new_n495_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n422_), .A2(KEYINPUT94), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n494_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n499_), .B1(new_n545_), .B2(new_n331_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT27), .B(new_n479_), .C1(new_n546_), .C2(new_n475_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n547_), .A2(KEYINPUT96), .A3(new_n536_), .A4(new_n537_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n531_), .A2(new_n542_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G227gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(G15gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT30), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n416_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT31), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT83), .B1(new_n432_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n555_), .B2(new_n432_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n554_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G71gat), .B(G99gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G43gat), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n560_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n549_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n547_), .A2(new_n536_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n563_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n486_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n565_), .A2(new_n568_), .A3(new_n529_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n572_));
  AND4_X1   g371(.A1(new_n206_), .A2(new_n204_), .A3(new_n211_), .A4(new_n209_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n224_), .A2(new_n225_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n219_), .A2(new_n205_), .A3(new_n214_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT15), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n291_), .B(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n572_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n227_), .A2(new_n295_), .A3(KEYINPUT73), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n228_), .A2(new_n291_), .A3(new_n230_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT34), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n583_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n589_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n581_), .A2(new_n584_), .A3(new_n582_), .A4(new_n590_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT77), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n592_), .A2(KEYINPUT77), .A3(new_n593_), .A4(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT36), .Z(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n595_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n325_), .A2(new_n571_), .A3(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n567_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n279_), .A2(new_n268_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT13), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n275_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT72), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n281_), .A2(KEYINPUT72), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n569_), .B1(new_n549_), .B2(new_n563_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n604_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT37), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n608_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n324_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR4_X1   g426(.A1(new_n619_), .A2(new_n309_), .A3(new_n620_), .A4(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n283_), .A3(new_n486_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n629_), .A2(KEYINPUT97), .A3(new_n611_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT97), .B1(new_n629_), .B2(new_n611_), .ZN(new_n631_));
  OAI221_X1 g430(.A(new_n610_), .B1(new_n611_), .B2(new_n629_), .C1(new_n630_), .C2(new_n631_), .ZN(G1324gat));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n284_), .B1(new_n633_), .B2(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(new_n565_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n609_), .B2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n638_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n635_), .A2(G8gat), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n639_), .A2(new_n640_), .B1(new_n628_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n642_), .B(new_n643_), .Z(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n609_), .B2(new_n563_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT41), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n628_), .A2(new_n551_), .A3(new_n566_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  OAI21_X1  g447(.A(G22gat), .B1(new_n609_), .B2(new_n530_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n628_), .A2(new_n651_), .A3(new_n529_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1327gat));
  NOR2_X1   g452(.A1(new_n620_), .A2(new_n309_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n281_), .A2(new_n608_), .A3(new_n626_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n486_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n281_), .A2(new_n309_), .A3(new_n626_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n625_), .B2(KEYINPUT100), .ZN(new_n660_));
  INV_X1    g459(.A(new_n604_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n662_), .A2(new_n598_), .B1(new_n606_), .B2(new_n595_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n622_), .B1(new_n663_), .B2(KEYINPUT37), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n660_), .B1(new_n571_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n620_), .A2(new_n668_), .A3(new_n625_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n659_), .B1(new_n665_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT44), .B(new_n659_), .C1(new_n665_), .C2(new_n669_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n486_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n658_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  NOR2_X1   g475(.A1(new_n635_), .A2(G36gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n657_), .A2(KEYINPUT103), .A3(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  INV_X1    g479(.A(new_n677_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n656_), .B2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n678_), .A2(new_n679_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n679_), .B1(new_n678_), .B2(new_n682_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n672_), .A2(new_n565_), .A3(new_n673_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G36gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G36gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT46), .B(new_n685_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1329gat));
  AOI21_X1  g493(.A(G43gat), .B1(new_n657_), .B2(new_n566_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n566_), .A2(G43gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n674_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1330gat));
  AOI21_X1  g498(.A(G50gat), .B1(new_n657_), .B2(new_n529_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n529_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n674_), .B2(new_n701_), .ZN(G1331gat));
  NOR4_X1   g501(.A1(new_n620_), .A2(new_n614_), .A3(new_n627_), .A4(new_n308_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n486_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n324_), .A2(new_n308_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR4_X1   g506(.A1(new_n618_), .A2(new_n620_), .A3(new_n663_), .A4(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n486_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n709_), .B2(new_n704_), .ZN(G1332gat));
  INV_X1    g509(.A(G64gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n708_), .B2(new_n565_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT48), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n703_), .A2(new_n711_), .A3(new_n565_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n708_), .B2(new_n566_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT105), .B(KEYINPUT49), .Z(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n703_), .A2(new_n716_), .A3(new_n566_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1334gat));
  INV_X1    g520(.A(G78gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n703_), .A2(new_n722_), .A3(new_n529_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n708_), .A2(new_n529_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(G78gat), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G78gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT107), .Z(G1335gat));
  NOR3_X1   g528(.A1(new_n618_), .A2(new_n608_), .A3(new_n626_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n620_), .A2(new_n308_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n486_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n626_), .A2(new_n308_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n281_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n665_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n669_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n486_), .A2(new_n202_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT108), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n734_), .B1(new_n739_), .B2(new_n741_), .ZN(G1336gat));
  INV_X1    g541(.A(new_n739_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G92gat), .B1(new_n743_), .B2(new_n635_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n732_), .A2(G92gat), .A3(new_n635_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n743_), .B2(new_n563_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n566_), .A2(new_n207_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n732_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n208_), .A3(new_n529_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n739_), .A2(new_n529_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G106gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT52), .B(new_n208_), .C1(new_n739_), .C2(new_n529_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n756_), .B(new_n758_), .ZN(G1339gat));
  NOR2_X1   g558(.A1(new_n565_), .A2(new_n529_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n486_), .A3(new_n566_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(KEYINPUT59), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n625_), .B(new_n706_), .C1(new_n276_), .C2(new_n280_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT111), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT54), .B1(new_n763_), .B2(new_n764_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n707_), .B1(new_n613_), .B2(new_n275_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n767_), .A2(KEYINPUT110), .A3(new_n768_), .A4(new_n625_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n765_), .A2(new_n766_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n765_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n268_), .A2(new_n308_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n251_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n245_), .B(KEYINPUT55), .C1(new_n249_), .C2(new_n250_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n245_), .A2(new_n246_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n256_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n278_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n278_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n773_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n292_), .A2(new_n293_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n293_), .B1(new_n297_), .B2(new_n291_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n296_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(new_n305_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n279_), .B2(new_n268_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n608_), .B1(new_n784_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT57), .B(new_n608_), .C1(new_n784_), .C2(new_n790_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n789_), .B1(new_n273_), .B2(new_n255_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n278_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n278_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT112), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n796_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT58), .B(new_n796_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n664_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n626_), .B1(new_n795_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n762_), .B1(new_n772_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n308_), .B2(KEYINPUT115), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(KEYINPUT115), .B2(new_n811_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n803_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n799_), .B2(KEYINPUT112), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n806_), .B1(new_n815_), .B2(new_n802_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n793_), .B(new_n794_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n324_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n765_), .A2(new_n769_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n766_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n765_), .A2(new_n766_), .A3(new_n769_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n761_), .B1(new_n820_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n810_), .B(new_n813_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n820_), .A2(new_n825_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n761_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n308_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n811_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT116), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n828_), .A2(new_n832_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1340gat));
  OAI211_X1 g636(.A(new_n619_), .B(new_n810_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n816_), .A2(new_n817_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n795_), .A3(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n842_), .A2(new_n324_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n843_), .B2(new_n761_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n619_), .A4(new_n810_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n839_), .A2(G120gat), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n614_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n826_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n826_), .B2(new_n626_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n853_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n844_), .A2(new_n810_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT119), .B(G127gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n626_), .A2(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(KEYINPUT120), .Z(new_n860_));
  AOI22_X1  g659(.A1(new_n854_), .A2(new_n855_), .B1(new_n857_), .B2(new_n860_), .ZN(G1342gat));
  OAI21_X1  g660(.A(G134gat), .B1(new_n856_), .B2(new_n625_), .ZN(new_n862_));
  INV_X1    g661(.A(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n826_), .A2(new_n863_), .A3(new_n663_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1343gat));
  NOR4_X1   g664(.A1(new_n565_), .A2(new_n530_), .A3(new_n567_), .A4(new_n566_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n829_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n309_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n437_), .ZN(G1344gat));
  INV_X1    g668(.A(new_n867_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n619_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT121), .B(G148gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n867_), .A2(new_n324_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OR3_X1    g675(.A1(new_n867_), .A2(G162gat), .A3(new_n608_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G162gat), .B1(new_n867_), .B2(new_n625_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n772_), .A2(new_n809_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n635_), .A2(new_n568_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n308_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT122), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n529_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n880_), .B1(new_n886_), .B2(G169gat), .ZN(new_n887_));
  AOI211_X1 g686(.A(KEYINPUT62), .B(new_n377_), .C1(new_n881_), .C2(new_n885_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n882_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n529_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n881_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n308_), .A2(new_n396_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT123), .Z(new_n893_));
  OAI22_X1  g692(.A1(new_n887_), .A2(new_n888_), .B1(new_n891_), .B2(new_n893_), .ZN(G1348gat));
  NAND3_X1  g693(.A1(new_n881_), .A2(new_n281_), .A3(new_n890_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n843_), .A2(new_n529_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n618_), .A2(new_n378_), .A3(new_n889_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n895_), .A2(new_n378_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  NAND2_X1  g697(.A1(new_n369_), .A2(new_n371_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n891_), .A2(new_n900_), .A3(new_n324_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n626_), .A3(new_n882_), .ZN(new_n902_));
  INV_X1    g701(.A(G183gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n891_), .B2(new_n625_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n663_), .A2(new_n370_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n891_), .B2(new_n906_), .ZN(G1351gat));
  NAND3_X1  g706(.A1(new_n565_), .A2(new_n563_), .A3(new_n537_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n843_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n308_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT124), .B(G197gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1352gat));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n619_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g713(.A(new_n324_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n909_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT125), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n916_), .A2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n918_), .B(KEYINPUT126), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n916_), .B2(new_n921_), .ZN(G1354gat));
  NOR2_X1   g721(.A1(new_n608_), .A2(G218gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n909_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n909_), .B2(new_n664_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT127), .B1(new_n925_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n843_), .A2(new_n625_), .A3(new_n908_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n924_), .B(new_n929_), .C1(new_n926_), .C2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n928_), .A2(new_n931_), .ZN(G1355gat));
endmodule


