//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n213_));
  OAI22_X1  g012(.A1(new_n212_), .A2(new_n213_), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT68), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n223_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n211_), .B1(new_n222_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n232_), .A2(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n221_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT65), .B1(new_n215_), .B2(new_n216_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT6), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n235_), .A2(new_n243_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n231_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT9), .B1(new_n224_), .B2(new_n225_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n247_), .B(KEYINPUT64), .C1(KEYINPUT9), .C2(new_n224_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT10), .B(G99gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n220_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n224_), .A2(new_n251_), .A3(KEYINPUT9), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n248_), .A2(new_n243_), .A3(new_n250_), .A4(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n210_), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n236_), .A2(new_n242_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n214_), .A2(new_n221_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n230_), .B(new_n245_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n222_), .A2(new_n230_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT8), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n209_), .A3(new_n253_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n255_), .A2(KEYINPUT12), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n253_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n210_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n255_), .A2(new_n262_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n268_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G120gat), .B(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT69), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n269_), .A2(new_n272_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n202_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(new_n279_), .A3(KEYINPUT13), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n284_), .A3(KEYINPUT70), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT71), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G232gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT34), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT35), .ZN(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G29gat), .B(G36gat), .ZN(new_n296_));
  INV_X1    g095(.A(G50gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G43gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n264_), .A2(new_n295_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n264_), .B2(new_n295_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n293_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n264_), .A2(new_n295_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n298_), .B(new_n299_), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n292_), .B(KEYINPUT35), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n311_));
  XOR2_X1   g110(.A(G134gat), .B(G162gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G190gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT77), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n310_), .A2(new_n319_), .A3(new_n311_), .A4(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n316_), .B(KEYINPUT36), .Z(new_n322_));
  NOR2_X1   g121(.A1(new_n310_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT37), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n321_), .A2(KEYINPUT37), .A3(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n209_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G1gat), .B(G8gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G15gat), .ZN(new_n335_));
  INV_X1    g134(.A(G22gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G15gat), .A2(G22gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G1gat), .A2(G8gat), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n337_), .A2(new_n338_), .B1(KEYINPUT14), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n334_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n331_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G183gat), .B(G211gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G127gat), .B(G155gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n343_), .B1(KEYINPUT17), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT80), .A3(KEYINPUT17), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n329_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n290_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT82), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n342_), .A2(new_n300_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n306_), .A2(new_n341_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n295_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G229gat), .A2(G233gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n300_), .A2(new_n294_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n341_), .B(new_n300_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(KEYINPUT83), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G113gat), .B(G141gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G169gat), .B(G197gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n365_), .A2(KEYINPUT83), .A3(new_n368_), .A4(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377_));
  INV_X1    g176(.A(G85gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT2), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G141gat), .A3(G148gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388_));
  NOR4_X1   g187(.A1(new_n388_), .A2(KEYINPUT88), .A3(G141gat), .A4(G148gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT89), .ZN(new_n394_));
  AND2_X1   g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n398_), .B(new_n387_), .C1(new_n389_), .C2(new_n392_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT1), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n390_), .B1(new_n395_), .B2(KEYINPUT1), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n383_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G127gat), .B(G134gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n400_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(KEYINPUT4), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT92), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n410_), .A2(KEYINPUT4), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n410_), .A2(new_n417_), .A3(KEYINPUT4), .A4(new_n411_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n410_), .A2(new_n414_), .A3(new_n411_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n382_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n419_), .A2(KEYINPUT93), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(KEYINPUT93), .ZN(new_n425_));
  AND4_X1   g224(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .A4(new_n382_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT24), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G169gat), .A2(G176gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n433_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n438_));
  AND2_X1   g237(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n438_), .A2(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G169gat), .ZN(new_n443_));
  INV_X1    g242(.A(G176gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT84), .A3(KEYINPUT24), .A4(new_n434_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT85), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G183gat), .A2(G190gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(KEYINPUT86), .A2(G183gat), .A3(G190gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT23), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n445_), .A2(KEYINPUT24), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n437_), .A2(new_n442_), .A3(new_n458_), .A4(new_n446_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n448_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT22), .B(G169gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n444_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n451_), .A2(KEYINPUT23), .A3(new_n452_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n449_), .A2(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G183gat), .A2(G190gat), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n434_), .B(new_n462_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT30), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(KEYINPUT30), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n409_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n408_), .A3(new_n469_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G43gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G227gat), .A2(G233gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n432_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n472_), .A2(new_n474_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n477_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n431_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n400_), .A2(new_n487_), .A3(new_n404_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(KEYINPUT28), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(KEYINPUT28), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n489_), .A2(new_n297_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n297_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G228gat), .A2(G233gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n487_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT21), .ZN(new_n499_));
  INV_X1    g298(.A(G197gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(G197gat), .B2(new_n274_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n274_), .A2(G197gat), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n499_), .B(new_n501_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G211gat), .B(G218gat), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n500_), .A2(G204gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT21), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT21), .A3(new_n506_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n495_), .B1(new_n498_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n495_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n510_), .A2(new_n512_), .ZN(new_n516_));
  NOR4_X1   g315(.A1(new_n496_), .A2(new_n497_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(G22gat), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(KEYINPUT90), .A3(new_n513_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n515_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n498_), .A2(new_n495_), .A3(new_n513_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n336_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n494_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n514_), .A2(new_n517_), .A3(G22gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n336_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n524_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n493_), .A3(new_n526_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n486_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G8gat), .B(G36gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G92gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT18), .B(G64gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G226gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT19), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n468_), .B2(new_n513_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n453_), .A2(new_n466_), .A3(new_n456_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n462_), .A2(new_n434_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n454_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n445_), .A2(KEYINPUT24), .A3(new_n434_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n442_), .A3(new_n547_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n544_), .A2(new_n545_), .B1(new_n548_), .B2(new_n465_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(new_n513_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n541_), .B1(new_n543_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n460_), .A2(new_n516_), .A3(new_n467_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n513_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(KEYINPUT20), .A3(new_n541_), .A4(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n539_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT27), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n516_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n559_), .A2(new_n542_), .A3(new_n550_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n555_), .B(new_n538_), .C1(new_n560_), .C2(new_n541_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n557_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(KEYINPUT96), .ZN(new_n563_));
  INV_X1    g362(.A(new_n541_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n549_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n549_), .A2(new_n565_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n516_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n568_), .B2(new_n543_), .ZN(new_n569_));
  AND4_X1   g368(.A1(KEYINPUT20), .A2(new_n553_), .A3(new_n564_), .A4(new_n554_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n538_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n539_), .C1(new_n552_), .C2(new_n556_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n563_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  AOI211_X1 g373(.A(KEYINPUT97), .B(new_n562_), .C1(new_n574_), .C2(KEYINPUT27), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(KEYINPUT27), .ZN(new_n577_));
  INV_X1    g376(.A(new_n562_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n534_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n533_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n493_), .B1(new_n532_), .B2(new_n526_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n562_), .B1(new_n574_), .B2(KEYINPUT27), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n486_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n428_), .B1(new_n580_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n486_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n555_), .B1(new_n560_), .B2(new_n541_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n590_), .B2(new_n538_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT32), .B(new_n539_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n591_), .B(new_n592_), .C1(new_n423_), .C2(new_n426_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n424_), .A2(new_n422_), .A3(new_n425_), .A4(new_n382_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n421_), .A2(new_n422_), .A3(new_n382_), .A4(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n557_), .A2(new_n561_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n410_), .A2(new_n415_), .A3(new_n411_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n381_), .A3(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .A4(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n588_), .B1(new_n593_), .B2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n359_), .B(new_n376_), .C1(new_n587_), .C2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n376_), .B1(new_n587_), .B2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT98), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n358_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(G1gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n428_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n587_), .A2(new_n604_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n321_), .A2(KEYINPUT99), .A3(new_n324_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT99), .B1(new_n321_), .B2(new_n324_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n355_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n289_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n376_), .A4(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n427_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n610_), .A2(new_n611_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n621_), .A3(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(new_n573_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n572_), .B1(new_n589_), .B2(new_n539_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n558_), .B1(new_n626_), .B2(new_n571_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT97), .B1(new_n627_), .B2(new_n562_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n584_), .A2(new_n576_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n620_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(G8gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT100), .B1(new_n631_), .B2(new_n632_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT39), .A3(new_n636_), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n633_), .A2(new_n634_), .A3(KEYINPUT39), .ZN(new_n638_));
  INV_X1    g437(.A(new_n630_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n608_), .A2(new_n632_), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n637_), .A2(new_n638_), .A3(KEYINPUT40), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  OAI21_X1  g444(.A(G15gat), .B1(new_n620_), .B2(new_n486_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT41), .Z(new_n647_));
  INV_X1    g446(.A(new_n486_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n608_), .A2(new_n335_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1326gat));
  XOR2_X1   g449(.A(new_n583_), .B(KEYINPUT101), .Z(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G22gat), .B1(new_n620_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n608_), .A2(new_n336_), .A3(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n289_), .B1(new_n607_), .B2(new_n605_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n616_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n618_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n661_), .B2(new_n427_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n327_), .A2(KEYINPUT103), .A3(new_n328_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT37), .B1(new_n321_), .B2(new_n324_), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n326_), .B(new_n323_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n587_), .B2(new_n604_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n593_), .A2(new_n603_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n588_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n529_), .A2(new_n486_), .A3(new_n533_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n584_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n630_), .B2(new_n534_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(new_n428_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n329_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n670_), .A2(KEYINPUT43), .B1(new_n677_), .B2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n287_), .A2(new_n355_), .A3(new_n376_), .A4(new_n288_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT102), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n663_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n683_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n678_), .B1(new_n677_), .B2(new_n669_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n613_), .A2(new_n679_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n685_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n684_), .A2(G29gat), .A3(new_n688_), .A4(new_n428_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n662_), .A2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n658_), .A2(new_n691_), .A3(new_n639_), .A4(new_n660_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT45), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n670_), .A2(KEYINPUT43), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n677_), .A2(new_n680_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n683_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n639_), .B1(new_n696_), .B2(KEYINPUT44), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n681_), .A2(new_n663_), .A3(new_n683_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G36gat), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT104), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n684_), .A2(new_n639_), .A3(new_n688_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(G36gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n693_), .A2(new_n700_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n701_), .A2(new_n702_), .A3(G36gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n702_), .B1(new_n701_), .B2(G36gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n712_), .A2(new_n705_), .A3(new_n706_), .A4(new_n693_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n709_), .A2(new_n713_), .ZN(G1329gat));
  NAND4_X1  g513(.A1(new_n684_), .A2(G43gat), .A3(new_n688_), .A4(new_n648_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n661_), .A2(new_n486_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G43gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g517(.A(new_n297_), .B1(new_n661_), .B2(new_n652_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n583_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n684_), .A2(G50gat), .A3(new_n688_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT106), .Z(G1331gat));
  INV_X1    g522(.A(new_n290_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n355_), .A2(new_n376_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n617_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n427_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n613_), .A2(new_n376_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT107), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n619_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n356_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n427_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n733_), .B2(new_n732_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n728_), .B1(new_n735_), .B2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n726_), .B2(new_n630_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT48), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n630_), .A2(G64gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n732_), .B2(new_n739_), .ZN(G1333gat));
  OR3_X1    g539(.A1(new_n732_), .A2(G71gat), .A3(new_n486_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n726_), .A2(new_n486_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G71gat), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n743_), .A2(KEYINPUT109), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(KEYINPUT109), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n741_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n726_), .B2(new_n652_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n732_), .A2(G78gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n652_), .ZN(G1335gat));
  NAND2_X1  g552(.A1(new_n694_), .A2(new_n695_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n376_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n619_), .A2(new_n618_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n757_), .A2(new_n378_), .A3(new_n427_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n660_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n730_), .A2(new_n290_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n428_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n761_), .B2(new_n378_), .ZN(G1336gat));
  AOI21_X1  g561(.A(G92gat), .B1(new_n760_), .B2(new_n639_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n757_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n639_), .A2(G92gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT110), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n764_), .B2(new_n766_), .ZN(G1337gat));
  NAND3_X1  g566(.A1(new_n760_), .A2(new_n249_), .A3(new_n648_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G99gat), .B1(new_n757_), .B2(new_n486_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g570(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(new_n583_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT52), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n220_), .A3(new_n583_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n772_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n776_), .B1(new_n773_), .B2(G106gat), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT52), .B(new_n220_), .C1(new_n764_), .C2(new_n583_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n779_), .B(new_n772_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n780_), .A2(new_n784_), .ZN(G1339gat));
  NOR2_X1   g584(.A1(new_n639_), .A2(new_n427_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n534_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT118), .ZN(new_n788_));
  INV_X1    g587(.A(new_n285_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n327_), .A2(new_n789_), .A3(new_n328_), .A4(new_n725_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT112), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT113), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n790_), .A2(KEYINPUT112), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n796_), .A3(new_n792_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n795_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT113), .B(KEYINPUT54), .C1(new_n790_), .C2(KEYINPUT112), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n804_));
  NAND3_X1  g603(.A1(new_n362_), .A2(new_n367_), .A3(new_n364_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n366_), .A2(new_n363_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n373_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n372_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n807_), .B(new_n808_), .C1(new_n283_), .C2(new_n279_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n269_), .A2(KEYINPUT114), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n271_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(KEYINPUT55), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n263_), .A2(new_n271_), .A3(new_n266_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n811_), .A2(new_n814_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n277_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n277_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n277_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n269_), .A2(new_n272_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n376_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n277_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(KEYINPUT115), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n809_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n804_), .B1(new_n829_), .B2(new_n616_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT117), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n616_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT57), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n807_), .A2(new_n808_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n822_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n834_), .B(new_n825_), .C1(new_n835_), .C2(new_n827_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n820_), .A2(new_n822_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n834_), .A4(new_n825_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n840_), .A3(new_n329_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n804_), .C1(new_n829_), .C2(new_n616_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n831_), .A2(new_n833_), .A3(new_n841_), .A4(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n355_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n788_), .B1(new_n803_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT119), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n798_), .A2(new_n802_), .B1(new_n844_), .B2(new_n355_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n849_), .B(KEYINPUT59), .C1(new_n850_), .C2(new_n788_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n830_), .A2(new_n853_), .A3(new_n841_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n833_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n830_), .B2(new_n841_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n355_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n803_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n788_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n847_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n858_), .A2(new_n862_), .A3(new_n847_), .A4(new_n859_), .ZN(new_n863_));
  INV_X1    g662(.A(G113gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n755_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n852_), .A2(new_n861_), .A3(new_n863_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n803_), .A2(new_n845_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n859_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n868_), .B2(new_n755_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n866_), .A2(new_n869_), .ZN(G1340gat));
  NAND4_X1  g669(.A1(new_n852_), .A2(new_n724_), .A3(new_n861_), .A4(new_n863_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT122), .B(G120gat), .Z(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n872_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n874_), .A2(KEYINPUT60), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT60), .B1(new_n289_), .B2(new_n874_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n868_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT123), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n873_), .A2(new_n878_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n355_), .A2(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n852_), .A2(new_n861_), .A3(new_n863_), .A4(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n868_), .B2(new_n355_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1342gat));
  INV_X1    g683(.A(new_n329_), .ZN(new_n885_));
  INV_X1    g684(.A(G134gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n852_), .A2(new_n861_), .A3(new_n863_), .A4(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n868_), .B2(new_n659_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n850_), .A2(new_n674_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n786_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n755_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT124), .B(G141gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  INV_X1    g694(.A(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n724_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g697(.A1(new_n892_), .A2(new_n355_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT61), .B(G155gat), .Z(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n896_), .B2(new_n616_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n669_), .A2(G162gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n896_), .B2(new_n903_), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n630_), .A2(new_n428_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n652_), .A2(new_n648_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n858_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n755_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n909_), .A2(new_n461_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n443_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT62), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n911_), .A2(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1348gat));
  NAND2_X1  g713(.A1(new_n867_), .A2(new_n720_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n905_), .A2(new_n648_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n915_), .A2(new_n444_), .A3(new_n290_), .A4(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n906_), .B1(new_n857_), .B2(new_n803_), .ZN(new_n918_));
  AOI21_X1  g717(.A(G176gat), .B1(new_n918_), .B2(new_n289_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1349gat));
  OR3_X1    g719(.A1(new_n915_), .A2(new_n355_), .A3(new_n916_), .ZN(new_n921_));
  INV_X1    g720(.A(G183gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n355_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n922_), .B1(new_n918_), .B2(new_n923_), .ZN(G1350gat));
  OAI211_X1 g723(.A(new_n918_), .B(new_n616_), .C1(new_n441_), .C2(new_n440_), .ZN(new_n925_));
  INV_X1    g724(.A(G190gat), .ZN(new_n926_));
  AOI211_X1 g725(.A(KEYINPUT125), .B(new_n926_), .C1(new_n918_), .C2(new_n329_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n858_), .A2(new_n329_), .A3(new_n907_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(G190gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n925_), .B1(new_n927_), .B2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT126), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n933_), .B(new_n925_), .C1(new_n927_), .C2(new_n930_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n891_), .A2(new_n905_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n755_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n500_), .ZN(G1352gat));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n290_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n274_), .ZN(G1353gat));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AND2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  NOR4_X1   g741(.A1(new_n936_), .A2(new_n355_), .A3(new_n941_), .A4(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n936_), .B2(new_n355_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  OAI211_X1 g745(.A(KEYINPUT127), .B(new_n941_), .C1(new_n936_), .C2(new_n355_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n943_), .B1(new_n946_), .B2(new_n947_), .ZN(G1354gat));
  INV_X1    g747(.A(new_n936_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n949_), .A2(G218gat), .A3(new_n329_), .ZN(new_n950_));
  AOI21_X1  g749(.A(G218gat), .B1(new_n949_), .B2(new_n616_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1355gat));
endmodule


