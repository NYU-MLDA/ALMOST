//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT82), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n207_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n208_), .A2(new_n209_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n216_), .B(KEYINPUT3), .Z(new_n220_));
  XOR2_X1   g019(.A(new_n218_), .B(KEYINPUT2), .Z(new_n221_));
  OAI211_X1 g020(.A(new_n211_), .B(new_n210_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G127gat), .A2(G134gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G120gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G127gat), .A2(G134gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  OAI21_X1  g028(.A(G120gat), .B1(new_n229_), .B2(new_n224_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT80), .B(G113gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n223_), .A2(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n232_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT90), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT90), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n242_), .A3(new_n235_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n241_), .A2(new_n243_), .A3(new_n219_), .A4(new_n222_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT91), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n204_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n236_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT4), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n203_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n202_), .A3(new_n248_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G1gat), .B(G29gat), .ZN(new_n254_));
  INV_X1    g053(.A(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n252_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n247_), .B1(new_n238_), .B2(new_n244_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n241_), .A2(new_n243_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n219_), .A2(new_n222_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT91), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n251_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n202_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n253_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n258_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT89), .ZN(new_n272_));
  INV_X1    g071(.A(G169gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT22), .B1(new_n273_), .B2(KEYINPUT79), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT79), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(G169gat), .ZN(new_n277_));
  INV_X1    g076(.A(G176gat), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT23), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(G183gat), .A3(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n281_), .A2(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n279_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n285_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n292_), .A2(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n288_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n281_), .A2(new_n283_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(KEYINPUT78), .A3(new_n303_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n301_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n290_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n310_), .A2(G197gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(G197gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT21), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(new_n318_), .A3(new_n314_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n309_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n286_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n287_), .B(KEYINPUT87), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n276_), .A2(new_n273_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT88), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n329_), .A3(new_n326_), .ZN(new_n330_));
  AOI21_X1  g129(.A(G176gat), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n319_), .B(new_n315_), .C1(new_n324_), .C2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT85), .B1(new_n297_), .B2(new_n300_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n304_), .ZN(new_n334_));
  AND2_X1   g133(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n337_));
  OAI22_X1  g136(.A1(new_n291_), .A2(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n273_), .A2(new_n278_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT24), .A3(new_n287_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n334_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT86), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n333_), .A2(new_n345_), .A3(new_n334_), .A4(new_n342_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n332_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n302_), .A2(KEYINPUT78), .A3(new_n303_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT78), .B1(new_n302_), .B2(new_n303_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n289_), .B1(new_n354_), .B2(new_n301_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n315_), .A2(new_n319_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n348_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n324_), .A2(new_n331_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n357_), .B1(new_n359_), .B2(new_n356_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n321_), .A2(new_n351_), .B1(new_n360_), .B2(new_n350_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G92gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT18), .B(G64gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  OAI21_X1  g164(.A(new_n272_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n332_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n338_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n339_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n345_), .B1(new_n370_), .B2(new_n334_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n346_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n367_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n350_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(KEYINPUT20), .A3(new_n374_), .A4(new_n321_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT20), .B1(new_n309_), .B2(new_n320_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n324_), .A2(new_n331_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n378_), .B2(new_n320_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n365_), .B(new_n375_), .C1(new_n379_), .C2(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n360_), .A2(new_n350_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n375_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n365_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT89), .A3(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n366_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT95), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n381_), .A2(KEYINPUT95), .A3(new_n365_), .A4(new_n375_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT27), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n368_), .A2(new_n369_), .A3(new_n304_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n332_), .C2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n321_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n377_), .A2(new_n356_), .A3(new_n343_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT93), .B1(new_n396_), .B2(KEYINPUT20), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n350_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n374_), .B(new_n357_), .C1(new_n359_), .C2(new_n356_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n392_), .B1(new_n400_), .B2(new_n383_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n391_), .A2(KEYINPUT96), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT96), .B1(new_n391_), .B2(new_n401_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n271_), .B(new_n387_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT28), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT84), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n408_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G22gat), .B(G50gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n356_), .B1(new_n223_), .B2(KEYINPUT29), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT83), .Z(new_n416_));
  OR2_X1    g215(.A1(new_n408_), .A2(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n410_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n412_), .A3(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n414_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n407_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n419_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n414_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n406_), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n309_), .A2(KEYINPUT30), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n309_), .A2(KEYINPUT30), .ZN(new_n429_));
  OAI21_X1  g228(.A(G43gat), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n309_), .A2(KEYINPUT30), .ZN(new_n431_));
  INV_X1    g230(.A(G43gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n309_), .A2(KEYINPUT30), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  AND3_X1   g237(.A1(new_n430_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT81), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n434_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n430_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n236_), .B(KEYINPUT31), .Z(new_n448_));
  NAND3_X1  g247(.A1(new_n441_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT81), .B(new_n450_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n422_), .A2(new_n427_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT98), .B1(new_n404_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT95), .B1(new_n361_), .B2(new_n365_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n390_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n401_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n391_), .A2(KEYINPUT96), .A3(new_n401_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n458_), .A2(new_n459_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT98), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n422_), .A2(new_n427_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n449_), .A2(new_n451_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n460_), .A2(new_n461_), .A3(new_n271_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n453_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n404_), .A2(new_n462_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n400_), .A2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n382_), .A2(new_n468_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n259_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n267_), .A2(new_n268_), .A3(new_n258_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n469_), .B(new_n470_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT94), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n366_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n250_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n248_), .B1(new_n477_), .B2(new_n247_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n251_), .B1(new_n478_), .B2(KEYINPUT4), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n476_), .B1(new_n479_), .B2(new_n203_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n246_), .A2(new_n203_), .A3(new_n248_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT92), .B(new_n202_), .C1(new_n249_), .C2(new_n251_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n480_), .A2(new_n258_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n260_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n472_), .A2(KEYINPUT33), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n475_), .A2(new_n483_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n462_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n270_), .A2(new_n489_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n474_), .A2(new_n487_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n467_), .A2(new_n491_), .A3(new_n463_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n466_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n255_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n503_), .A2(new_n510_), .A3(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT66), .B(KEYINPUT9), .ZN(new_n513_));
  INV_X1    g312(.A(new_n506_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT67), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT9), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT66), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n516_), .B(new_n506_), .C1(new_n518_), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(KEYINPUT9), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n515_), .A2(new_n505_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n500_), .A2(new_n501_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT10), .B(G99gat), .Z(new_n525_));
  AOI21_X1  g324(.A(new_n524_), .B1(new_n525_), .B2(new_n496_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n512_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT68), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n512_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G57gat), .ZN(new_n532_));
  INV_X1    g331(.A(G64gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT11), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G57gat), .A2(G64gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538_));
  INV_X1    g337(.A(G71gat), .ZN(new_n539_));
  INV_X1    g338(.A(G78gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT69), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n535_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT69), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n537_), .A2(new_n545_), .A3(new_n538_), .A4(new_n541_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n529_), .A2(new_n531_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n512_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n530_), .B1(new_n512_), .B2(new_n527_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n553_), .A2(new_n554_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT70), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n512_), .A2(new_n527_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n512_), .B2(new_n527_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT12), .B(new_n549_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n552_), .A2(new_n555_), .A3(new_n558_), .A4(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n555_), .A2(new_n550_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n558_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G120gat), .B(G148gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(G204gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT5), .B(G176gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n571_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(KEYINPUT13), .A3(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G15gat), .B(G22gat), .Z(new_n579_));
  NAND2_X1  g378(.A1(G1gat), .A2(G8gat), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(KEYINPUT14), .B2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT76), .ZN(new_n582_));
  XOR2_X1   g381(.A(G1gat), .B(G8gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G43gat), .B(G50gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G29gat), .B(G36gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT15), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n582_), .A2(new_n583_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n587_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n582_), .A2(new_n583_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n584_), .A2(new_n587_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n594_), .A3(KEYINPUT77), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT77), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n584_), .A2(new_n598_), .A3(new_n587_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(new_n600_), .B2(new_n590_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n601_), .B(new_n604_), .Z(new_n605_));
  NOR2_X1   g404(.A1(new_n578_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n493_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n588_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n592_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n608_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n611_), .A2(new_n613_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n618_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT74), .ZN(new_n622_));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT36), .ZN(new_n626_));
  INV_X1    g425(.A(new_n621_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT36), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT73), .Z(new_n630_));
  AOI22_X1  g429(.A1(new_n622_), .A2(new_n626_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n630_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n621_), .A2(new_n626_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n631_), .A2(new_n632_), .B1(KEYINPUT37), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n549_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(new_n584_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G127gat), .B(G155gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT16), .B(G183gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(new_n642_), .Z(new_n643_));
  INV_X1    g442(.A(KEYINPUT17), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n639_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n645_), .B2(new_n639_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n636_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n607_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G1gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n270_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n631_), .A2(new_n649_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n607_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n271_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n658_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(G8gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n460_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n655_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n607_), .A2(new_n666_), .A3(new_n660_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(G8gat), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT102), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n670_), .A2(new_n675_), .A3(G8gat), .A4(new_n671_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n673_), .A2(new_n674_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n667_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n667_), .B(KEYINPUT40), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  OAI21_X1  g482(.A(G15gat), .B1(new_n661_), .B2(new_n463_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT41), .Z(new_n685_));
  INV_X1    g484(.A(G15gat), .ZN(new_n686_));
  INV_X1    g485(.A(new_n463_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n653_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1326gat));
  OAI21_X1  g488(.A(G22gat), .B1(new_n661_), .B2(new_n488_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT42), .ZN(new_n691_));
  INV_X1    g490(.A(G22gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n653_), .A2(new_n692_), .A3(new_n462_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n622_), .A2(new_n626_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n633_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n648_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n607_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n270_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n466_), .A2(new_n701_), .A3(new_n492_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n466_), .B2(new_n492_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n700_), .B1(new_n704_), .B2(new_n636_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n493_), .A2(new_n700_), .A3(new_n636_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n493_), .A2(KEYINPUT104), .A3(new_n700_), .A4(new_n636_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n606_), .B(new_n649_), .C1(new_n705_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n270_), .A2(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n699_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n666_), .A3(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n698_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n460_), .A2(KEYINPUT105), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n460_), .A2(KEYINPUT105), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n720_), .A2(G36gat), .A3(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n719_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n719_), .A2(KEYINPUT46), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  NAND4_X1  g532(.A1(new_n713_), .A2(new_n714_), .A3(G43gat), .A4(new_n687_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT107), .B(G43gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n720_), .B2(new_n463_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g537(.A1(new_n713_), .A2(new_n462_), .A3(new_n714_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT108), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(KEYINPUT108), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(G50gat), .A3(new_n741_), .ZN(new_n742_));
  OR3_X1    g541(.A1(new_n720_), .A2(G50gat), .A3(new_n488_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n493_), .A2(new_n605_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT109), .Z(new_n746_));
  INV_X1    g545(.A(new_n578_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n270_), .A3(new_n650_), .ZN(new_n749_));
  AND4_X1   g548(.A1(new_n605_), .A2(new_n493_), .A3(new_n578_), .A4(new_n660_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n271_), .A2(new_n532_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n749_), .A2(new_n532_), .B1(new_n750_), .B2(new_n751_), .ZN(G1332gat));
  AOI21_X1  g551(.A(new_n533_), .B1(new_n750_), .B2(new_n724_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n748_), .A2(new_n650_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n724_), .A2(new_n533_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(G1333gat));
  AOI21_X1  g557(.A(new_n539_), .B1(new_n750_), .B2(new_n687_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT49), .Z(new_n760_));
  NAND2_X1  g559(.A1(new_n687_), .A2(new_n539_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT111), .Z(G1334gat));
  AOI21_X1  g562(.A(new_n540_), .B1(new_n750_), .B2(new_n462_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT50), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n462_), .A2(new_n540_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n756_), .B2(new_n766_), .ZN(G1335gat));
  AND2_X1   g566(.A1(new_n748_), .A2(new_n697_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n270_), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n705_), .A2(new_n710_), .A3(KEYINPUT112), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n601_), .B(new_n604_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n747_), .A2(new_n771_), .A3(new_n648_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n705_), .B2(new_n710_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n270_), .A2(G85gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT113), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n769_), .B1(new_n774_), .B2(new_n776_), .ZN(G1336gat));
  AOI21_X1  g576(.A(G92gat), .B1(new_n768_), .B2(new_n666_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n725_), .A2(new_n504_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n774_), .B2(new_n779_), .ZN(G1337gat));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT51), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n781_), .A2(KEYINPUT51), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G99gat), .B1(new_n784_), .B2(new_n463_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n768_), .A2(new_n525_), .A3(new_n687_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n782_), .B(new_n783_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  AND4_X1   g586(.A1(new_n781_), .A2(new_n785_), .A3(KEYINPUT51), .A4(new_n786_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1338gat));
  OAI211_X1 g588(.A(new_n462_), .B(new_n772_), .C1(new_n705_), .C2(new_n710_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(KEYINPUT52), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n768_), .A2(new_n496_), .A3(new_n462_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n792_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .A4(new_n800_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n601_), .A2(new_n604_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n589_), .A2(new_n594_), .ZN(new_n806_));
  MUX2_X1   g605(.A(new_n806_), .B(new_n600_), .S(new_n590_), .Z(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n604_), .B2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n574_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n562_), .A2(new_n555_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n553_), .A2(new_n554_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT12), .B1(new_n811_), .B2(new_n549_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n565_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT55), .A3(new_n563_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n810_), .A2(new_n812_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n558_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n571_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT118), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n814_), .A2(new_n821_), .A3(new_n817_), .A4(new_n571_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT119), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n818_), .A2(new_n820_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n819_), .A2(new_n826_), .A3(new_n820_), .A4(new_n822_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n771_), .A2(new_n572_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n809_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT120), .B1(new_n830_), .B2(new_n631_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT57), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n818_), .B(new_n820_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n572_), .A3(new_n808_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n635_), .A2(KEYINPUT37), .ZN(new_n837_));
  INV_X1    g636(.A(new_n632_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n696_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT121), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n834_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT58), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n636_), .B(new_n843_), .C1(KEYINPUT58), .C2(new_n841_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(new_n842_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT120), .B(new_n846_), .C1(new_n830_), .C2(new_n631_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n832_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n605_), .A2(new_n577_), .A3(new_n576_), .A4(new_n648_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n839_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(KEYINPUT54), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT54), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n848_), .A2(new_n649_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n855_), .A2(new_n271_), .A3(new_n666_), .A4(new_n452_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n771_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n605_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g660(.A(new_n226_), .B1(new_n747_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT122), .B1(new_n226_), .B2(KEYINPUT60), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n856_), .B(new_n864_), .C1(new_n865_), .C2(new_n862_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n747_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n226_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n856_), .B2(new_n648_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n649_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g670(.A(G134gat), .B1(new_n856_), .B2(new_n631_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n839_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g673(.A1(new_n848_), .A2(new_n649_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n853_), .A2(new_n854_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n488_), .A2(new_n687_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n724_), .A2(new_n271_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n878_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n855_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(KEYINPUT123), .A3(new_n879_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n771_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n578_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT124), .B(G148gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1345gat));
  NAND2_X1  g690(.A1(new_n886_), .A2(new_n648_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  AOI21_X1  g693(.A(KEYINPUT123), .B1(new_n884_), .B2(new_n879_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n879_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n855_), .A2(new_n881_), .A3(new_n883_), .A4(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(G162gat), .B(new_n636_), .C1(new_n895_), .C2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n696_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT125), .B1(new_n900_), .B2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n631_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n899_), .B1(new_n901_), .B2(new_n905_), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n855_), .A2(new_n452_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n725_), .A2(new_n270_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n771_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G169gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT127), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n912_), .A3(G169gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n914_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n910_), .A2(KEYINPUT127), .A3(new_n916_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n328_), .A2(new_n330_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n909_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n915_), .A2(new_n917_), .A3(new_n919_), .ZN(G1348gat));
  NAND2_X1  g719(.A1(new_n907_), .A2(new_n908_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n747_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n278_), .ZN(G1349gat));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n649_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n291_), .B2(new_n335_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n284_), .B2(new_n924_), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n921_), .B2(new_n839_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n631_), .B1(new_n337_), .B2(new_n336_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n921_), .B2(new_n928_), .ZN(G1351gat));
  NAND2_X1  g728(.A1(new_n884_), .A2(new_n908_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n771_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n930_), .A2(new_n747_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n310_), .ZN(G1353gat));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n930_), .A2(new_n649_), .A3(new_n936_), .A4(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n931_), .A2(new_n648_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n936_), .ZN(G1354gat));
  AND3_X1   g739(.A1(new_n931_), .A2(G218gat), .A3(new_n636_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G218gat), .B1(new_n931_), .B2(new_n631_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1355gat));
endmodule


