//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT79), .B(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n210_), .B1(new_n216_), .B2(KEYINPUT80), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT80), .B2(new_n216_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n205_), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n220_), .B(KEYINPUT81), .Z(new_n221_));
  INV_X1    g020(.A(G183gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n212_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n203_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n208_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G227gat), .A2(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(G71gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G99gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT82), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT30), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT31), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n236_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT1), .Z(new_n247_));
  NOR2_X1   g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT83), .ZN(new_n249_));
  AOI211_X1 g048(.A(new_n243_), .B(new_n245_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n244_), .B(KEYINPUT2), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252_));
  OAI22_X1  g051(.A1(new_n252_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(KEYINPUT84), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT85), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n251_), .A2(new_n258_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n249_), .A2(new_n246_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n250_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G22gat), .B(G50gat), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT29), .B(new_n270_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n272_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G228gat), .A2(G233gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n283_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n284_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT90), .Z(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n262_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n264_), .A2(KEYINPUT29), .A3(new_n265_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n290_), .B(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(new_n281_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n282_), .A2(new_n294_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n280_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n279_), .A2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n299_), .A2(new_n301_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n279_), .A2(new_n304_), .A3(KEYINPUT91), .A4(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n264_), .A2(new_n235_), .A3(new_n265_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n262_), .A2(new_n311_), .A3(new_n234_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n262_), .A2(new_n234_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT94), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT4), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n310_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n317_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT33), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n327_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT33), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT26), .B(G190gat), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n211_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(new_n203_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n208_), .A3(new_n220_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n344_), .B2(new_n290_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n226_), .A2(new_n297_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT92), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT92), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n226_), .A2(new_n297_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n336_), .B1(new_n344_), .B2(new_n290_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n226_), .B2(new_n297_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n352_), .A2(new_n335_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G8gat), .B(G36gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n331_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n314_), .A2(new_n312_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n319_), .B1(new_n368_), .B2(new_n310_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n320_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n317_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT95), .B(new_n331_), .C1(new_n315_), .C2(new_n317_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n367_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n330_), .A2(new_n333_), .A3(new_n364_), .A4(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n350_), .A2(new_n353_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n347_), .A2(new_n349_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n291_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT20), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n335_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n352_), .A2(new_n335_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n376_), .B1(new_n383_), .B2(new_n375_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n321_), .A2(new_n331_), .A3(new_n322_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n332_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n309_), .B1(new_n374_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n321_), .A2(new_n331_), .A3(new_n322_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n328_), .A2(KEYINPUT96), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT96), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n385_), .B2(new_n332_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n383_), .A2(new_n359_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n392_), .A2(new_n394_), .B1(new_n363_), .B2(new_n393_), .ZN(new_n395_));
  AND4_X1   g194(.A1(new_n389_), .A2(new_n309_), .A3(new_n391_), .A4(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n242_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n309_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n395_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n389_), .A3(new_n241_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G232gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT34), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT35), .ZN(new_n406_));
  XOR2_X1   g205(.A(G29gat), .B(G36gat), .Z(new_n407_));
  XOR2_X1   g206(.A(G43gat), .B(G50gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT15), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT8), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT7), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT65), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT6), .ZN(new_n418_));
  AND2_X1   g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G99gat), .A2(G106gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n417_), .A2(KEYINPUT6), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n415_), .A2(KEYINPUT65), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G85gat), .B(G92gat), .Z(new_n426_));
  AOI21_X1  g225(.A(new_n412_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n412_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n414_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n419_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n424_), .A2(KEYINPUT66), .A3(new_n420_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n431_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n430_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI211_X1 g238(.A(KEYINPUT67), .B(new_n431_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n428_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n433_), .A2(new_n434_), .A3(new_n432_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT66), .B1(new_n424_), .B2(new_n420_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT64), .B(G92gat), .Z(new_n445_));
  INV_X1    g244(.A(KEYINPUT9), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(G85gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n426_), .A2(KEYINPUT9), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT10), .B(G99gat), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n447_), .B(new_n448_), .C1(G106gat), .C2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n411_), .B1(new_n441_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n406_), .B1(new_n453_), .B2(KEYINPUT71), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n441_), .A2(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n410_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n441_), .A2(new_n452_), .A3(new_n457_), .A4(new_n409_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n414_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n429_), .B1(new_n460_), .B2(KEYINPUT67), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n437_), .A2(new_n438_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n451_), .B1(new_n463_), .B2(new_n428_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n464_), .B2(new_n409_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n454_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n405_), .A2(KEYINPUT35), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n464_), .B2(new_n411_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n469_), .B2(new_n406_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n409_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT70), .B1(new_n455_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n458_), .A3(new_n456_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n466_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT74), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n466_), .B(KEYINPUT74), .C1(new_n470_), .C2(new_n473_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G190gat), .B(G218gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT72), .ZN(new_n479_));
  XOR2_X1   g278(.A(G134gat), .B(G162gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT36), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n476_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n481_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(KEYINPUT36), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n403_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G120gat), .B(G148gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  XOR2_X1   g294(.A(G71gat), .B(G78gat), .Z(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n427_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n451_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n441_), .A2(new_n452_), .A3(new_n500_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(KEYINPUT12), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT12), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n455_), .A2(new_n506_), .A3(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n493_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n509_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n493_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT69), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n513_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n510_), .A2(new_n512_), .A3(new_n493_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n516_), .B1(new_n515_), .B2(new_n511_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT69), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT13), .B1(new_n519_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n518_), .B1(new_n513_), .B2(new_n517_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT13), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(KEYINPUT69), .A3(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529_));
  INV_X1    g328(.A(G1gat), .ZN(new_n530_));
  INV_X1    g329(.A(G8gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G8gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n409_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT78), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(KEYINPUT78), .A3(new_n409_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n535_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n538_), .A2(new_n539_), .B1(new_n471_), .B2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n410_), .A2(new_n540_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G169gat), .B(G197gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  OR3_X1    g349(.A1(new_n544_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n528_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n500_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT75), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n535_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT77), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n566_));
  OR3_X1    g365(.A1(new_n558_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n554_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n488_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT97), .B1(new_n488_), .B2(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n391_), .A2(new_n389_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n403_), .A2(new_n554_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n474_), .A2(KEYINPUT73), .A3(new_n485_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n466_), .B(new_n482_), .C1(new_n470_), .C2(new_n473_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT73), .B1(new_n474_), .B2(new_n485_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n483_), .A2(new_n586_), .A3(new_n486_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n569_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n580_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n530_), .A3(new_n577_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n579_), .A2(new_n592_), .ZN(G1324gat));
  NOR3_X1   g392(.A1(new_n488_), .A2(new_n395_), .A3(new_n570_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n531_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n568_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n395_), .A2(G8gat), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n403_), .A2(new_n554_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT98), .Z(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(new_n594_), .B2(new_n531_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n596_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT40), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n596_), .A2(new_n600_), .A3(new_n605_), .A4(new_n601_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1325gat));
  NAND2_X1  g408(.A1(new_n575_), .A2(new_n241_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G15gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(G15gat), .A3(new_n612_), .ZN(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n590_), .A2(new_n616_), .A3(new_n241_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n614_), .A2(new_n615_), .A3(KEYINPUT102), .A4(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  NOR2_X1   g421(.A1(new_n398_), .A2(G22gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT103), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n590_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n576_), .B2(new_n398_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT42), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT42), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(G1327gat));
  NOR3_X1   g428(.A1(new_n580_), .A2(new_n487_), .A3(new_n569_), .ZN(new_n630_));
  INV_X1    g429(.A(G29gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n577_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n588_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n364_), .B(new_n373_), .C1(new_n332_), .C2(KEYINPUT33), .ZN(new_n635_));
  INV_X1    g434(.A(new_n333_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n386_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n398_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n309_), .A2(new_n391_), .A3(new_n395_), .A4(new_n389_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n241_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n633_), .B(new_n634_), .C1(new_n640_), .C2(new_n401_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n588_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n554_), .A2(new_n568_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n644_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n578_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n632_), .B1(new_n651_), .B2(new_n631_), .ZN(G1328gat));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n395_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n630_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT45), .ZN(new_n656_));
  INV_X1    g455(.A(new_n650_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n644_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n654_), .A4(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n649_), .A2(new_n650_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n658_), .B1(new_n662_), .B2(new_n654_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n656_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OAI221_X1 g466(.A(new_n656_), .B1(new_n665_), .B2(KEYINPUT46), .C1(new_n661_), .C2(new_n663_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  INV_X1    g468(.A(G43gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n630_), .A2(new_n670_), .A3(new_n241_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n649_), .A2(new_n650_), .A3(new_n242_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n670_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g473(.A(G50gat), .B1(new_n630_), .B2(new_n309_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n309_), .A2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n662_), .B2(new_n676_), .ZN(G1331gat));
  INV_X1    g476(.A(new_n528_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n553_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n403_), .A2(new_n597_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(G57gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n577_), .ZN(new_n683_));
  NOR4_X1   g482(.A1(new_n488_), .A2(new_n568_), .A3(new_n679_), .A4(new_n678_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(new_n577_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n685_), .B2(new_n682_), .ZN(G1332gat));
  INV_X1    g485(.A(G64gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n684_), .B2(new_n654_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT48), .Z(new_n689_));
  NOR2_X1   g488(.A1(new_n395_), .A2(G64gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT108), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n681_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1333gat));
  AOI21_X1  g492(.A(new_n228_), .B1(new_n684_), .B2(new_n241_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT49), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n228_), .A3(new_n241_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1334gat));
  INV_X1    g496(.A(G78gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n684_), .B2(new_n309_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n681_), .A2(new_n698_), .A3(new_n309_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1335gat));
  INV_X1    g502(.A(new_n487_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n403_), .A2(new_n704_), .A3(new_n568_), .A4(new_n680_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT110), .Z(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n577_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n644_), .A2(new_n568_), .A3(new_n680_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n577_), .A2(G85gat), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT111), .Z(new_n710_));
  AOI21_X1  g509(.A(new_n707_), .B1(new_n708_), .B2(new_n710_), .ZN(G1336gat));
  AOI21_X1  g510(.A(G92gat), .B1(new_n706_), .B2(new_n654_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n654_), .A2(new_n445_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n708_), .B2(new_n713_), .ZN(G1337gat));
  INV_X1    g513(.A(new_n449_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n706_), .A2(new_n241_), .A3(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n708_), .A2(new_n241_), .ZN(new_n717_));
  INV_X1    g516(.A(G99gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n719_), .B(new_n720_), .Z(G1338gat));
  INV_X1    g520(.A(G106gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(new_n722_), .A3(new_n309_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n708_), .A2(new_n309_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G106gat), .ZN(new_n726_));
  AOI211_X1 g525(.A(KEYINPUT52), .B(new_n722_), .C1(new_n708_), .C2(new_n309_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n723_), .B(new_n729_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1339gat));
  NAND3_X1  g532(.A1(new_n523_), .A2(new_n553_), .A3(new_n527_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n589_), .A2(KEYINPUT54), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT54), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n523_), .A2(new_n553_), .A3(new_n527_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n597_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n545_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n550_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n740_), .B(new_n741_), .C1(new_n542_), .C2(new_n541_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n552_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n524_), .A2(new_n526_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n524_), .A2(new_n745_), .A3(KEYINPUT115), .A4(new_n526_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n505_), .A2(new_n514_), .A3(new_n507_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n510_), .A2(KEYINPUT55), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n493_), .B1(new_n515_), .B2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n753_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n679_), .B(new_n520_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n748_), .A2(new_n749_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n487_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(KEYINPUT57), .A3(new_n487_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n756_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n754_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n745_), .A2(new_n520_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT58), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n588_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n765_), .A3(KEYINPUT58), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n761_), .A2(new_n762_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n739_), .B1(new_n770_), .B2(new_n568_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n399_), .A2(new_n578_), .A3(new_n242_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n679_), .ZN(new_n775_));
  INV_X1    g574(.A(G113gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n759_), .A2(new_n760_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n569_), .B1(new_n782_), .B2(new_n762_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT59), .B(new_n772_), .C1(new_n783_), .C2(new_n739_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n553_), .A2(new_n776_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n778_), .A2(new_n779_), .B1(new_n785_), .B2(new_n786_), .ZN(G1340gat));
  NOR2_X1   g586(.A1(new_n678_), .A2(KEYINPUT60), .ZN(new_n788_));
  INV_X1    g587(.A(G120gat), .ZN(new_n789_));
  MUX2_X1   g588(.A(KEYINPUT60), .B(new_n788_), .S(new_n789_), .Z(new_n790_));
  NAND2_X1  g589(.A1(new_n774_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n774_), .A2(KEYINPUT117), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n678_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  OAI21_X1  g596(.A(G120gat), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT118), .B(new_n678_), .C1(new_n781_), .C2(new_n784_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n795_), .B(KEYINPUT119), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1341gat));
  AOI21_X1  g603(.A(G127gat), .B1(new_n774_), .B2(new_n569_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n569_), .A2(G127gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT120), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n785_), .B2(new_n807_), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n774_), .A2(new_n809_), .A3(new_n704_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n588_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n809_), .ZN(G1343gat));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n398_), .A2(new_n654_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n577_), .A3(new_n242_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n771_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n815_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT121), .B(new_n817_), .C1(new_n783_), .C2(new_n739_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n679_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n528_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT122), .B(G148gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1345gat));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n819_), .B2(new_n569_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n819_), .A2(new_n825_), .A3(new_n569_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1346gat));
  INV_X1    g631(.A(new_n819_), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n833_), .A2(G162gat), .A3(new_n487_), .ZN(new_n834_));
  OAI21_X1  g633(.A(G162gat), .B1(new_n833_), .B2(new_n588_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n400_), .A2(new_n395_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT124), .Z(new_n838_));
  NOR3_X1   g637(.A1(new_n771_), .A2(new_n309_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n204_), .B1(new_n839_), .B2(new_n679_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n840_), .A2(KEYINPUT62), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n219_), .A3(new_n679_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(KEYINPUT62), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(G1348gat));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n528_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n569_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n847_), .A2(KEYINPUT125), .A3(new_n211_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT125), .B1(new_n847_), .B2(new_n211_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n222_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(G1350gat));
  NAND2_X1  g650(.A1(new_n839_), .A2(new_n633_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G190gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n839_), .A2(new_n339_), .A3(new_n704_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1351gat));
  INV_X1    g654(.A(new_n771_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n577_), .A2(new_n398_), .A3(new_n395_), .A4(new_n241_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n553_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT126), .B(G197gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1352gat));
  INV_X1    g660(.A(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n528_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n569_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  AND2_X1   g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n865_), .B2(new_n866_), .ZN(G1354gat));
  OAI21_X1  g668(.A(G218gat), .B1(new_n858_), .B2(new_n588_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n487_), .A2(G218gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n858_), .B2(new_n871_), .ZN(G1355gat));
endmodule


