//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n204_), .A2(new_n206_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT84), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n208_), .A3(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n215_), .A3(KEYINPUT85), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(new_n202_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n219_), .B(KEYINPUT31), .Z(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT86), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(KEYINPUT86), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G227gat), .A2(G233gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n223_), .B(G15gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT30), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G71gat), .B(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G43gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n225_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT23), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(G183gat), .A3(G190gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n233_), .A3(KEYINPUT83), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n235_), .A3(KEYINPUT23), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT78), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT78), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n234_), .B(new_n236_), .C1(new_n241_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247_));
  OR3_X1    g046(.A1(new_n247_), .A2(KEYINPUT82), .A3(G169gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT82), .B1(new_n247_), .B2(G169gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(G176gat), .B1(new_n247_), .B2(G169gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n245_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n231_), .A2(new_n233_), .ZN(new_n253_));
  INV_X1    g052(.A(G169gat), .ZN(new_n254_));
  INV_X1    g053(.A(G176gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT24), .A3(new_n246_), .ZN(new_n257_));
  OR3_X1    g056(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(KEYINPUT81), .B2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n261_), .A2(KEYINPUT81), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n238_), .A2(new_n240_), .A3(KEYINPUT25), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n242_), .A2(KEYINPUT26), .A3(new_n243_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n237_), .B2(KEYINPUT25), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n267_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n259_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n252_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n229_), .B(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n221_), .A2(new_n222_), .A3(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n222_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280_));
  XOR2_X1   g079(.A(G155gat), .B(G162gat), .Z(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT3), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT89), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT88), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n288_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n289_), .B1(new_n288_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n281_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n283_), .A2(new_n284_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(KEYINPUT1), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n302_), .A2(KEYINPUT1), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n301_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n297_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n219_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n211_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n215_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n297_), .B(new_n310_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n280_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n297_), .A2(new_n310_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(KEYINPUT4), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n316_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n315_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n317_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n320_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n315_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT4), .B1(new_n330_), .B2(new_n318_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n317_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n319_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n327_), .B1(new_n334_), .B2(new_n322_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n279_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT94), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n297_), .A2(new_n310_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT28), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n297_), .A2(new_n310_), .A3(new_n345_), .A4(new_n342_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G22gat), .B(G50gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n344_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n341_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n347_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n339_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n344_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n342_), .B1(new_n297_), .B2(new_n310_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358_));
  INV_X1    g157(.A(G211gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(G218gat), .ZN(new_n360_));
  INV_X1    g159(.A(G218gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(G211gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT21), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT21), .ZN(new_n367_));
  AND2_X1   g166(.A1(G197gat), .A2(G204gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G197gat), .A2(G204gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n368_), .A2(new_n369_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n372_), .B(KEYINPUT21), .C1(new_n362_), .C2(new_n360_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n371_), .A2(KEYINPUT91), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT91), .B1(new_n371_), .B2(new_n373_), .ZN(new_n375_));
  INV_X1    g174(.A(G228gat), .ZN(new_n376_));
  INV_X1    g175(.A(G233gat), .ZN(new_n377_));
  OAI22_X1  g176(.A1(new_n374_), .A2(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT92), .B1(new_n357_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n376_), .A2(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n371_), .A2(new_n373_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT91), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n288_), .A2(new_n294_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT89), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n288_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n309_), .B1(new_n390_), .B2(new_n281_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n385_), .B(new_n386_), .C1(new_n391_), .C2(new_n342_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n379_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n381_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n380_), .B1(new_n357_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT93), .B(new_n380_), .C1(new_n357_), .C2(new_n394_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n351_), .A2(new_n356_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n245_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n269_), .A2(new_n271_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(new_n264_), .A3(new_n267_), .A4(new_n265_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n259_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n383_), .A2(new_n405_), .A3(new_n409_), .A4(new_n384_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n253_), .B1(G183gat), .B2(G190gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n246_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n255_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT25), .B(G183gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n261_), .A2(G190gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n260_), .A2(KEYINPUT26), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT95), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n260_), .A2(KEYINPUT26), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n261_), .A2(G190gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n417_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n234_), .A2(new_n257_), .A3(new_n236_), .A4(new_n258_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n415_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n381_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n410_), .A2(KEYINPUT20), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT19), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT18), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n426_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n424_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n423_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n416_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n437_), .A2(new_n440_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT96), .A3(new_n394_), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n252_), .A2(new_n273_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT96), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n427_), .B2(new_n381_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n431_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .A4(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n432_), .A2(new_n436_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n436_), .B1(new_n432_), .B2(new_n448_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n404_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  INV_X1    g251(.A(new_n436_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n431_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n410_), .A2(KEYINPUT20), .A3(new_n428_), .A4(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n446_), .B1(new_n441_), .B2(new_n394_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(new_n443_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n432_), .A2(new_n436_), .A3(new_n448_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT27), .A3(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n451_), .A2(new_n452_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n452_), .B1(new_n451_), .B2(new_n461_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n402_), .B(new_n403_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n432_), .A2(new_n448_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n453_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT27), .B1(new_n467_), .B2(new_n460_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n459_), .A2(KEYINPUT27), .A3(new_n460_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT99), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n451_), .A2(new_n452_), .A3(new_n461_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n403_), .B1(new_n472_), .B2(new_n402_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n338_), .B1(new_n465_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n401_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n351_), .A2(new_n356_), .A3(new_n399_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n468_), .A2(new_n469_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n477_), .A2(new_n336_), .A3(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n328_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT33), .B(new_n328_), .C1(new_n320_), .C2(new_n323_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n327_), .B1(new_n321_), .B2(new_n317_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n317_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT97), .B(new_n327_), .C1(new_n321_), .C2(new_n317_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n449_), .A2(new_n450_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n482_), .A2(new_n483_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n432_), .A2(new_n492_), .A3(new_n448_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n456_), .A2(new_n458_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n466_), .B2(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n329_), .B2(new_n335_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n477_), .B1(new_n491_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n278_), .B1(new_n479_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n474_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G85gat), .B(G92gat), .Z(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n504_), .A2(KEYINPUT9), .ZN(new_n517_));
  INV_X1    g316(.A(G85gat), .ZN(new_n518_));
  INV_X1    g317(.A(G92gat), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT9), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n510_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT10), .B(G99gat), .Z(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT64), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT64), .B1(new_n522_), .B2(new_n523_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n517_), .B(new_n521_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n511_), .A2(new_n512_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n528_), .B1(KEYINPUT8), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT66), .B1(new_n516_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n525_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n521_), .A2(new_n517_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n515_), .A2(new_n513_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n514_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(KEYINPUT8), .A3(new_n529_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT12), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n531_), .A2(new_n538_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n516_), .A2(new_n530_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n545_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n546_), .B1(new_n516_), .B2(new_n530_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n534_), .A2(new_n536_), .A3(new_n545_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n551_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT67), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n557_), .A2(new_n560_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n564_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(KEYINPUT13), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT13), .B1(new_n567_), .B2(new_n569_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT75), .ZN(new_n574_));
  XOR2_X1   g373(.A(G15gat), .B(G22gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT70), .B(G1gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(G8gat), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n575_), .B1(new_n577_), .B2(KEYINPUT14), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G1gat), .B(G8gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n578_), .B(KEYINPUT71), .ZN(new_n583_));
  INV_X1    g382(.A(new_n581_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G29gat), .B(G36gat), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT68), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G43gat), .B(G50gat), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n582_), .A2(new_n585_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n574_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n592_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n583_), .A2(new_n584_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n580_), .A2(new_n581_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n582_), .A2(new_n585_), .A3(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(KEYINPUT75), .A3(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n595_), .A2(new_n601_), .A3(G229gat), .A4(G233gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT76), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n592_), .B(KEYINPUT15), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n582_), .A2(new_n585_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n599_), .B(new_n604_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT77), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n602_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(KEYINPUT77), .A3(new_n612_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n503_), .A2(new_n573_), .A3(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n620_));
  NAND2_X1  g419(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT36), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT34), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT35), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT15), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n592_), .B(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n552_), .A2(new_n596_), .B1(new_n630_), .B2(new_n629_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n632_), .A3(new_n636_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n626_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n635_), .A2(new_n632_), .A3(new_n636_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n641_), .A2(new_n637_), .A3(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n620_), .B(new_n621_), .C1(new_n640_), .C2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n642_), .A3(new_n639_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n625_), .B1(new_n641_), .B2(new_n637_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(KEYINPUT69), .A4(KEYINPUT37), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G127gat), .B(G155gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT16), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT74), .Z(new_n656_));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n545_), .B(new_n657_), .Z(new_n658_));
  XNOR2_X1  g457(.A(new_n606_), .B(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT72), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n660_), .B2(new_n659_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n653_), .B(KEYINPUT17), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n649_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n619_), .A2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n667_), .A2(new_n336_), .A3(new_n576_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT38), .Z(new_n669_));
  NOR2_X1   g468(.A1(new_n640_), .A2(new_n644_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n665_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n619_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n336_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(G1324gat));
  INV_X1    g473(.A(G8gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n672_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n472_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT101), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT39), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(KEYINPUT101), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n678_), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n619_), .A2(new_n675_), .A3(new_n677_), .A4(new_n666_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n682_), .A2(KEYINPUT40), .A3(new_n683_), .A4(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n680_), .A2(new_n681_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n684_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(new_n689_), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n672_), .B2(new_n278_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT41), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n667_), .A2(G15gat), .A3(new_n278_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n672_), .B2(new_n402_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n402_), .A2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n667_), .B2(new_n698_), .ZN(G1327gat));
  OAI21_X1  g498(.A(new_n402_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT100), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n337_), .B1(new_n701_), .B2(new_n464_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n483_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n335_), .A2(KEYINPUT33), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n500_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n402_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n477_), .A2(new_n336_), .A3(new_n478_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n279_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n649_), .B1(new_n702_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n649_), .C1(new_n702_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n573_), .A2(new_n618_), .A3(new_n665_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n717_), .B(new_n714_), .C1(new_n710_), .C2(new_n712_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n720_));
  INV_X1    g519(.A(new_n336_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n670_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n665_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n619_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n336_), .A2(G29gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT104), .Z(new_n730_));
  OAI22_X1  g529(.A1(new_n723_), .A2(new_n724_), .B1(new_n728_), .B2(new_n730_), .ZN(G1328gat));
  AOI21_X1  g530(.A(new_n711_), .B1(new_n503_), .B2(new_n649_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n712_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n715_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n717_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n715_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n677_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n728_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n677_), .A2(KEYINPUT106), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n677_), .A2(KEYINPUT106), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n739_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n728_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n738_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT105), .B1(new_n737_), .B2(G36gat), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT107), .B(KEYINPUT46), .C1(new_n750_), .C2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n716_), .A2(new_n718_), .A3(new_n472_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n743_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n738_), .A3(new_n749_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT46), .B1(new_n757_), .B2(KEYINPUT107), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n753_), .A2(new_n758_), .ZN(G1329gat));
  NOR3_X1   g558(.A1(new_n716_), .A2(new_n718_), .A3(new_n278_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n227_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n279_), .A2(new_n227_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n728_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g564(.A(G50gat), .B1(new_n739_), .B2(new_n477_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n477_), .A2(G50gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n719_), .B2(new_n767_), .ZN(G1331gat));
  NAND2_X1  g567(.A1(new_n567_), .A2(new_n569_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT13), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n570_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n666_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT108), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n618_), .B1(new_n474_), .B2(new_n502_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT109), .Z(new_n777_));
  INV_X1    g576(.A(G57gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n721_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n772_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n780_), .A2(new_n665_), .A3(new_n670_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G57gat), .B1(new_n782_), .B2(new_n336_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n783_), .ZN(G1332gat));
  INV_X1    g583(.A(G64gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n777_), .A2(new_n785_), .A3(new_n742_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n781_), .B2(new_n742_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT48), .Z(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1333gat));
  INV_X1    g588(.A(G71gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n781_), .B2(new_n279_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT49), .Z(new_n792_));
  NAND2_X1  g591(.A1(new_n279_), .A2(new_n790_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT110), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n777_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(G1334gat));
  INV_X1    g595(.A(G78gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n781_), .B2(new_n477_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT111), .Z(new_n799_));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n800_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n777_), .A2(new_n797_), .A3(new_n477_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(G1335gat));
  NOR3_X1   g603(.A1(new_n780_), .A2(new_n726_), .A3(new_n725_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n518_), .A3(new_n721_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n616_), .A2(new_n617_), .ZN(new_n807_));
  AND4_X1   g606(.A1(new_n772_), .A2(new_n713_), .A3(new_n807_), .A4(new_n665_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n721_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n809_), .B2(new_n518_), .ZN(G1336gat));
  NAND3_X1  g609(.A1(new_n805_), .A2(new_n519_), .A3(new_n677_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n808_), .A2(new_n742_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n519_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT112), .Z(G1337gat));
  INV_X1    g613(.A(G99gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n808_), .B2(new_n279_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n805_), .A2(new_n522_), .A3(new_n279_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n816_), .A2(new_n817_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n818_));
  NAND2_X1  g617(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n805_), .A2(new_n523_), .A3(new_n477_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n808_), .A2(new_n477_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(G106gat), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT52), .B(new_n523_), .C1(new_n808_), .C2(new_n477_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n771_), .A2(new_n570_), .A3(new_n807_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n645_), .A2(new_n648_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n726_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n573_), .A2(new_n666_), .A3(KEYINPUT114), .A4(new_n807_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(KEYINPUT54), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n828_), .B(new_n835_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n616_), .A2(new_n567_), .A3(new_n617_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n549_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n549_), .A2(new_n558_), .A3(new_n556_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n839_), .A2(KEYINPUT55), .B1(new_n551_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT115), .B1(new_n839_), .B2(KEYINPUT55), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n557_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n842_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n564_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n838_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n595_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n599_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n852_), .B(new_n612_), .C1(new_n853_), .C2(new_n604_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(new_n615_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n769_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n725_), .B1(new_n851_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n564_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n618_), .B(new_n567_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n856_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(KEYINPUT57), .A3(new_n725_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n862_), .A2(new_n861_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n861_), .A2(new_n867_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n567_), .A2(new_n855_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT117), .B(new_n866_), .C1(new_n868_), .C2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n649_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n870_), .B1(new_n867_), .B2(new_n861_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n849_), .A2(KEYINPUT116), .A3(new_n850_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n866_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n860_), .B(new_n865_), .C1(new_n874_), .C2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n837_), .B1(new_n880_), .B2(new_n665_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n701_), .A2(new_n464_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n721_), .A3(new_n279_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(G113gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n618_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n883_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n830_), .B1(new_n878_), .B2(new_n866_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n866_), .B2(new_n878_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n864_), .B2(new_n725_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n859_), .B(new_n670_), .C1(new_n863_), .C2(new_n856_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n726_), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT59), .B(new_n889_), .C1(new_n895_), .C2(new_n837_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n807_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n886_), .B1(new_n897_), .B2(new_n885_), .ZN(G1340gat));
  INV_X1    g697(.A(G120gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n884_), .B(new_n900_), .C1(KEYINPUT60), .C2(new_n899_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n573_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903_));
  OAI21_X1  g702(.A(G120gat), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  AOI211_X1 g703(.A(KEYINPUT118), .B(new_n573_), .C1(new_n888_), .C2(new_n896_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n901_), .B1(new_n904_), .B2(new_n905_), .ZN(G1341gat));
  AOI21_X1  g705(.A(G127gat), .B1(new_n884_), .B2(new_n726_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n888_), .A2(new_n896_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n665_), .A2(KEYINPUT119), .ZN(new_n909_));
  MUX2_X1   g708(.A(KEYINPUT119), .B(new_n909_), .S(G127gat), .Z(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(new_n908_), .B2(new_n910_), .ZN(G1342gat));
  NAND3_X1  g710(.A1(new_n884_), .A2(new_n203_), .A3(new_n670_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n830_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n203_), .ZN(G1343gat));
  INV_X1    g713(.A(new_n742_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n721_), .A3(new_n477_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n278_), .B(new_n917_), .C1(new_n895_), .C2(new_n837_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n807_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n283_), .ZN(G1344gat));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n918_), .B2(new_n573_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n881_), .A2(new_n279_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n922_), .A2(new_n923_), .A3(new_n772_), .A4(new_n917_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT120), .B(G148gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n921_), .A2(new_n924_), .A3(new_n926_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1345gat));
  NOR2_X1   g729(.A1(new_n918_), .A2(new_n665_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n931_), .B(new_n932_), .Z(G1346gat));
  INV_X1    g732(.A(G162gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n918_), .A2(new_n934_), .A3(new_n830_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n918_), .B2(new_n725_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT122), .B(new_n934_), .C1(new_n918_), .C2(new_n725_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1347gat));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n881_), .A2(new_n477_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n915_), .A2(new_n337_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n618_), .ZN(new_n944_));
  XOR2_X1   g743(.A(new_n944_), .B(KEYINPUT123), .Z(new_n945_));
  NAND2_X1  g744(.A1(new_n942_), .A2(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n941_), .B1(new_n946_), .B2(G169gat), .ZN(new_n947_));
  AOI211_X1 g746(.A(KEYINPUT62), .B(new_n254_), .C1(new_n942_), .C2(new_n945_), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n402_), .B(new_n943_), .C1(new_n895_), .C2(new_n837_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n618_), .A2(new_n413_), .ZN(new_n950_));
  OAI22_X1  g749(.A1(new_n947_), .A2(new_n948_), .B1(new_n949_), .B2(new_n950_), .ZN(G1348gat));
  NOR2_X1   g750(.A1(new_n949_), .A2(new_n573_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(new_n255_), .ZN(G1349gat));
  NOR2_X1   g752(.A1(new_n949_), .A2(new_n665_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n241_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n417_), .B2(new_n954_), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n949_), .B2(new_n830_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n725_), .B1(new_n424_), .B2(new_n420_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n942_), .A2(new_n943_), .A3(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(KEYINPUT124), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n957_), .A2(new_n962_), .A3(new_n959_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(G1351gat));
  NAND3_X1  g763(.A1(new_n742_), .A2(new_n336_), .A3(new_n477_), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n881_), .A2(new_n279_), .A3(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n618_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n772_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g769(.A(new_n665_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(KEYINPUT125), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n973_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n972_), .A2(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n966_), .A2(new_n975_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n973_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n977_));
  XOR2_X1   g776(.A(new_n976_), .B(new_n977_), .Z(G1354gat));
  NAND2_X1  g777(.A1(new_n966_), .A2(new_n670_), .ZN(new_n979_));
  XNOR2_X1  g778(.A(KEYINPUT127), .B(G218gat), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n830_), .A2(new_n980_), .ZN(new_n981_));
  AOI22_X1  g780(.A1(new_n979_), .A2(new_n980_), .B1(new_n966_), .B2(new_n981_), .ZN(G1355gat));
endmodule


