//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT99), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G64gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT81), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G169gat), .A3(G176gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT22), .B(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n216_), .B2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(KEYINPUT23), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G197gat), .B(G204gat), .Z(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n232_), .B(KEYINPUT21), .C1(KEYINPUT90), .C2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(KEYINPUT21), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT21), .B1(new_n233_), .B2(KEYINPUT90), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n231_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n223_), .ZN(new_n238_));
  NOR3_X1   g037(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n241_), .B2(new_n210_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n222_), .A2(new_n219_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G183gat), .ZN(new_n245_));
  INV_X1    g044(.A(G183gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT25), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(G190gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT26), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n245_), .A2(new_n247_), .A3(new_n249_), .A4(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n238_), .A2(new_n242_), .A3(new_n243_), .A4(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n230_), .A2(new_n234_), .A3(new_n237_), .A4(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(KEYINPUT80), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT26), .B(G190gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(KEYINPUT80), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n246_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(KEYINPUT79), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n241_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n239_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT23), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n225_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n262_), .B(new_n263_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n219_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n243_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n269_), .A2(new_n227_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272_));
  OR3_X1    g071(.A1(new_n272_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n273_));
  INV_X1    g072(.A(G176gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(G169gat), .B1(new_n272_), .B2(KEYINPUT83), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n214_), .ZN(new_n277_));
  OAI22_X1  g076(.A1(new_n261_), .A2(new_n268_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n237_), .A2(new_n234_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT92), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT19), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n254_), .A2(new_n280_), .A3(KEYINPUT20), .A4(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n227_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n253_), .B1(new_n286_), .B2(new_n217_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n285_), .B1(new_n287_), .B2(new_n279_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n239_), .B1(new_n214_), .B2(new_n241_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(new_n226_), .C1(new_n260_), .C2(new_n257_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n238_), .A2(new_n228_), .A3(new_n243_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n214_), .A3(new_n276_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n290_), .A2(new_n292_), .A3(new_n234_), .A4(new_n237_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n283_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n284_), .B1(new_n294_), .B2(KEYINPUT93), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  AOI211_X1 g095(.A(new_n296_), .B(new_n283_), .C1(new_n288_), .C2(new_n293_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n209_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(KEYINPUT94), .B(new_n209_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n294_), .A2(KEYINPUT93), .ZN(new_n302_));
  INV_X1    g101(.A(new_n297_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n284_), .A4(new_n208_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT98), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(KEYINPUT98), .A3(new_n306_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n288_), .A2(new_n283_), .A3(new_n293_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n254_), .A2(KEYINPUT20), .A3(new_n280_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n283_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n306_), .B1(new_n313_), .B2(new_n209_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n309_), .A2(new_n310_), .B1(new_n304_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G155gat), .B(G162gat), .Z(new_n316_));
  OR3_X1    g115(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n317_), .B(new_n318_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n316_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  OR2_X1    g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n323_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n279_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G228gat), .A3(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n279_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT91), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n323_), .A2(new_n329_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n341_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n333_), .A2(new_n335_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n336_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n338_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n339_), .A2(new_n348_), .A3(new_n338_), .A4(new_n345_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT96), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G113gat), .B(G120gat), .Z(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT87), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G113gat), .B(G120gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(G127gat), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(KEYINPUT87), .ZN(new_n362_));
  INV_X1    g161(.A(G127gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n359_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n361_), .A2(G134gat), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(G134gat), .B1(new_n361_), .B2(new_n365_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n340_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G134gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(G134gat), .A3(new_n365_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n330_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(KEYINPUT4), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n330_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n355_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT0), .ZN(new_n381_));
  INV_X1    g180(.A(G57gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n354_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n387_));
  OR3_X1    g186(.A1(new_n379_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n379_), .B2(new_n387_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n352_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n305_), .A2(KEYINPUT95), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n300_), .A2(new_n393_), .A3(new_n301_), .A4(new_n304_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n366_), .A2(new_n367_), .A3(new_n340_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT97), .B1(new_n395_), .B2(new_n376_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n368_), .A2(new_n397_), .A3(new_n374_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n354_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n375_), .A2(new_n355_), .A3(new_n378_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n399_), .A2(new_n385_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n389_), .A2(KEYINPUT33), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(new_n386_), .C1(new_n379_), .C2(new_n387_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n392_), .A2(new_n394_), .A3(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n208_), .A2(KEYINPUT32), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n313_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n302_), .A2(new_n303_), .A3(new_n284_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n390_), .B(new_n408_), .C1(new_n409_), .C2(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n315_), .A2(new_n391_), .B1(new_n411_), .B2(new_n352_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n278_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n417_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n366_), .A2(new_n367_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT31), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n426_), .A2(KEYINPUT86), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n426_), .B2(KEYINPUT86), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n423_), .A2(new_n424_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n424_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n428_), .A2(new_n429_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n422_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n203_), .B1(new_n412_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n314_), .A2(new_n304_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n305_), .A2(KEYINPUT98), .A3(new_n306_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT98), .B1(new_n305_), .B2(new_n306_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n391_), .B(new_n437_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n352_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT99), .B(new_n434_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n352_), .B(new_n437_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n434_), .A2(new_n445_), .A3(new_n390_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n436_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  INV_X1    g248(.A(G99gat), .ZN(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n452_), .A2(new_n455_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n384_), .A2(new_n207_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT66), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n464_), .A3(new_n461_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(KEYINPUT8), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n455_), .A2(new_n456_), .ZN(new_n469_));
  XOR2_X1   g268(.A(KEYINPUT10), .B(G99gat), .Z(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n451_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n459_), .A3(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n467_), .A2(new_n468_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n466_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT67), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(KEYINPUT11), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(KEYINPUT12), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n466_), .A2(new_n477_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n479_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n479_), .A2(new_n486_), .A3(new_n488_), .A4(KEYINPUT68), .ZN(new_n492_));
  INV_X1    g291(.A(new_n484_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n478_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n485_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT64), .ZN(new_n497_));
  INV_X1    g296(.A(new_n478_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(new_n484_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n491_), .A2(new_n492_), .A3(new_n495_), .A4(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n494_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n497_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n505_));
  XNOR2_X1  g304(.A(G120gat), .B(G148gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n500_), .A2(new_n503_), .A3(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT13), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(KEYINPUT13), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G8gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT74), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT75), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(G15gat), .A2(G22gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G15gat), .A2(G22gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G1gat), .A2(G8gat), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n524_), .A2(new_n525_), .B1(KEYINPUT14), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n520_), .A2(new_n521_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n520_), .A2(new_n521_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G29gat), .B(G36gat), .Z(new_n534_));
  XOR2_X1   g333(.A(G43gat), .B(G50gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT15), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT78), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT78), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n529_), .A2(new_n537_), .A3(new_n540_), .A4(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n532_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n536_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n536_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n529_), .A2(new_n549_), .A3(new_n532_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n542_), .A2(new_n545_), .B1(new_n551_), .B2(new_n544_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  INV_X1    g352(.A(G169gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G197gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n552_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n517_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n533_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n566_), .A2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n484_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n493_), .A3(new_n568_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT17), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n565_), .B1(new_n574_), .B2(new_n563_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT77), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n575_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n558_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT36), .Z(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT34), .Z(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n479_), .A2(new_n537_), .A3(new_n488_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT70), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(new_n587_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT71), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n478_), .B2(new_n549_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT72), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n589_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n590_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n598_), .A2(new_n588_), .A3(new_n595_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n584_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT73), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n583_), .A2(KEYINPUT36), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n597_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n604_), .B(new_n584_), .C1(new_n597_), .C2(new_n599_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n448_), .A2(new_n580_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n202_), .B1(new_n608_), .B2(new_n390_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n603_), .A2(new_n600_), .A3(KEYINPUT37), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n448_), .A2(new_n580_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n202_), .A3(new_n390_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n609_), .B1(new_n610_), .B2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n610_), .B2(new_n617_), .ZN(G1324gat));
  INV_X1    g418(.A(G8gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n315_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n448_), .A2(new_n621_), .A3(new_n580_), .A4(new_n606_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n622_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(G1325gat));
  OR3_X1    g431(.A1(new_n615_), .A2(G15gat), .A3(new_n434_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n608_), .A2(new_n435_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(new_n634_), .B2(G15gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(G1326gat));
  OR3_X1    g436(.A1(new_n615_), .A2(G22gat), .A3(new_n352_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G22gat), .B1(new_n607_), .B2(new_n352_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT42), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT42), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(G1327gat));
  AND3_X1   g441(.A1(new_n436_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n606_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n558_), .A2(new_n578_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n390_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n645_), .B(KEYINPUT102), .Z(new_n649_));
  OAI21_X1  g448(.A(new_n434_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n446_), .B1(new_n650_), .B2(new_n203_), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT43), .B(new_n614_), .C1(new_n651_), .C2(new_n444_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  INV_X1    g452(.A(new_n606_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n611_), .B1(new_n654_), .B2(KEYINPUT37), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n448_), .B2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n649_), .B(KEYINPUT44), .C1(new_n652_), .C2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(G29gat), .A3(new_n390_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n652_), .A2(new_n656_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n645_), .B(KEYINPUT102), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n648_), .B1(new_n658_), .B2(new_n662_), .ZN(G1328gat));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n643_), .B2(new_n614_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n448_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n661_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n315_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n669_), .B2(new_n662_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n315_), .A2(G36gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n647_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT45), .B1(new_n646_), .B2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n664_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n668_), .A2(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n657_), .A2(new_n621_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G36gat), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n673_), .A2(new_n675_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(KEYINPUT46), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n682_), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n657_), .A2(G43gat), .A3(new_n435_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n646_), .A2(new_n434_), .ZN(new_n685_));
  OAI22_X1  g484(.A1(new_n684_), .A2(new_n678_), .B1(G43gat), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n647_), .B2(new_n442_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n657_), .A2(G50gat), .A3(new_n442_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g489(.A(new_n517_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n578_), .ZN(new_n692_));
  NOR4_X1   g491(.A1(new_n643_), .A2(new_n557_), .A3(new_n654_), .A4(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n382_), .B1(new_n693_), .B2(new_n390_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n655_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT103), .Z(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(new_n643_), .A3(new_n557_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n390_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(G57gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n694_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT104), .ZN(G1332gat));
  INV_X1    g500(.A(G64gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n702_), .A3(new_n621_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n693_), .A2(new_n621_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G64gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT105), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n707_), .A3(G64gat), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n706_), .A2(KEYINPUT48), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT48), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n703_), .B1(new_n709_), .B2(new_n710_), .ZN(G1333gat));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n693_), .B2(new_n435_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT49), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n697_), .A2(new_n712_), .A3(new_n435_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1334gat));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n693_), .B2(new_n442_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT50), .Z(new_n719_));
  NAND3_X1  g518(.A1(new_n697_), .A2(new_n717_), .A3(new_n442_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1335gat));
  NOR3_X1   g520(.A1(new_n517_), .A2(new_n578_), .A3(new_n557_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n722_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT106), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n722_), .C1(new_n652_), .C2(new_n656_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n698_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n644_), .A2(new_n722_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n390_), .A2(new_n384_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n727_), .A2(new_n384_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  OAI21_X1  g529(.A(new_n207_), .B1(new_n728_), .B2(new_n315_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT107), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n724_), .A2(new_n726_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n315_), .A2(new_n207_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1337gat));
  NAND4_X1  g534(.A1(new_n644_), .A2(new_n435_), .A3(new_n470_), .A4(new_n722_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n434_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n450_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT51), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n738_), .B(new_n742_), .C1(new_n739_), .C2(new_n450_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1338gat));
  NAND4_X1  g543(.A1(new_n644_), .A2(new_n451_), .A3(new_n442_), .A4(new_n722_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n442_), .B(new_n722_), .C1(new_n652_), .C2(new_n656_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n745_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1339gat));
  NAND3_X1  g553(.A1(new_n542_), .A2(new_n548_), .A3(new_n544_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n556_), .B1(new_n551_), .B2(new_n543_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n552_), .A2(new_n556_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n512_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT111), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n760_), .A3(new_n512_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  OR3_X1    g562(.A1(new_n500_), .A2(KEYINPUT109), .A3(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n491_), .A2(new_n501_), .A3(new_n492_), .A4(new_n495_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n763_), .A2(new_n500_), .B1(new_n765_), .B2(new_n497_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT109), .B1(new_n500_), .B2(new_n763_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n510_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n510_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n762_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n762_), .B(KEYINPUT58), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n655_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n557_), .A2(new_n512_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n770_), .B2(new_n769_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n513_), .A2(new_n757_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n654_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(KEYINPUT57), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n579_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n557_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n614_), .A2(new_n517_), .A3(new_n785_), .A4(new_n578_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT54), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n435_), .A2(new_n390_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n445_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n792_), .B2(new_n791_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n788_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n791_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n780_), .B2(KEYINPUT57), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n768_), .A2(new_n510_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n510_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n776_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n779_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n606_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT110), .A3(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n798_), .A2(new_n807_), .A3(new_n781_), .A4(new_n775_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n579_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n796_), .B1(new_n809_), .B2(new_n787_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n795_), .B1(new_n810_), .B2(new_n789_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n785_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n810_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n785_), .A2(G113gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(G1340gat));
  OAI211_X1 g614(.A(new_n795_), .B(new_n691_), .C1(new_n810_), .C2(new_n789_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G120gat), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n517_), .A2(G120gat), .ZN(new_n818_));
  MUX2_X1   g617(.A(new_n818_), .B(G120gat), .S(KEYINPUT60), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n817_), .A2(KEYINPUT113), .A3(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1341gat));
  AOI21_X1  g624(.A(G127gat), .B1(new_n810_), .B2(new_n578_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n811_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n578_), .A2(G127gat), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT114), .Z(new_n829_));
  AOI21_X1  g628(.A(new_n826_), .B1(new_n827_), .B2(new_n829_), .ZN(G1342gat));
  NAND2_X1  g629(.A1(new_n655_), .A2(G134gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT115), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n811_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(G134gat), .B1(new_n810_), .B2(new_n654_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT116), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n834_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n836_), .B(new_n837_), .C1(new_n811_), .C2(new_n832_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1343gat));
  NAND4_X1  g638(.A1(new_n315_), .A2(new_n434_), .A3(new_n442_), .A4(new_n390_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n809_), .B2(new_n787_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n557_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n691_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT117), .B(G148gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT118), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n844_), .B(new_n846_), .ZN(G1345gat));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n578_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  INV_X1    g649(.A(G162gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n841_), .A2(new_n851_), .A3(new_n654_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n841_), .A2(new_n655_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1347gat));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n315_), .A2(new_n434_), .A3(new_n390_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n352_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n554_), .B1(new_n858_), .B2(new_n557_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT62), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n215_), .A3(new_n557_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n859_), .B2(KEYINPUT62), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n855_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n859_), .A2(KEYINPUT62), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT119), .A3(new_n860_), .A4(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1348gat));
  AOI21_X1  g666(.A(G176gat), .B1(new_n858_), .B2(new_n691_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n442_), .B1(new_n809_), .B2(new_n787_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n856_), .A2(new_n691_), .A3(G176gat), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n869_), .A2(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  INV_X1    g672(.A(new_n858_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n259_), .A3(new_n579_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n578_), .A3(new_n856_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G183gat), .B1(new_n876_), .B2(new_n877_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(G1350gat));
  NOR2_X1   g679(.A1(new_n874_), .A2(new_n614_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n250_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n654_), .A2(new_n256_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT122), .Z(new_n884_));
  NOR2_X1   g683(.A1(new_n874_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT123), .B1(new_n882_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  OAI221_X1 g686(.A(new_n887_), .B1(new_n874_), .B2(new_n884_), .C1(new_n881_), .C2(new_n250_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1351gat));
  NAND2_X1  g688(.A1(new_n809_), .A2(new_n787_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n621_), .A2(new_n434_), .A3(new_n391_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n557_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT124), .B(G204gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n691_), .ZN(new_n897_));
  MUX2_X1   g696(.A(new_n895_), .B(new_n896_), .S(new_n897_), .Z(G1353gat));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n579_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n892_), .A2(new_n899_), .A3(new_n900_), .A4(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n890_), .A2(new_n891_), .A3(new_n901_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(KEYINPUT125), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT126), .B1(new_n904_), .B2(KEYINPUT125), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n902_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n902_), .B2(new_n906_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1354gat));
  NAND2_X1  g708(.A1(new_n892_), .A2(new_n654_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT127), .B(G218gat), .Z(new_n911_));
  NOR2_X1   g710(.A1(new_n614_), .A2(new_n911_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n892_), .B2(new_n912_), .ZN(G1355gat));
endmodule


