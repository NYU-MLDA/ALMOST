//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT80), .B(G183gat), .Z(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT23), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n207_), .A2(KEYINPUT83), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(KEYINPUT83), .B2(new_n207_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n204_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n212_), .C1(new_n219_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n209_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G183gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(G190gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(KEYINPUT25), .B2(new_n208_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n223_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n214_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G197gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G204gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT88), .ZN(new_n237_));
  INV_X1    g036(.A(G204gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G197gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT87), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT21), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(new_n239_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n202_), .B1(new_n234_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT19), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n219_), .B1(KEYINPUT93), .B2(new_n222_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n222_), .A2(KEYINPUT93), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n211_), .B(KEYINPUT23), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n221_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT92), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT25), .B(G183gat), .Z(new_n264_));
  OAI211_X1 g063(.A(new_n259_), .B(new_n261_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n212_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n206_), .A3(new_n205_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n253_), .B(new_n256_), .C1(new_n252_), .C2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n252_), .A2(new_n268_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n214_), .A2(new_n248_), .A3(new_n233_), .A4(new_n251_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT20), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n255_), .B(KEYINPUT91), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT95), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n269_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n280_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT98), .B1(new_n265_), .B2(new_n267_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(new_n252_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(new_n268_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n256_), .B1(new_n292_), .B2(new_n253_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n272_), .A2(new_n273_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n288_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n284_), .A2(new_n285_), .B1(new_n287_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297_));
  INV_X1    g096(.A(G43gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n214_), .B2(new_n233_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G134gat), .Z(new_n303_));
  XOR2_X1   g102(.A(G113gat), .B(G120gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n214_), .A2(new_n233_), .A3(new_n300_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n305_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n306_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(new_n301_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G227gat), .A2(G233gat), .ZN(new_n312_));
  INV_X1    g111(.A(G15gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT30), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT31), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n307_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326_));
  INV_X1    g125(.A(G141gat), .ZN(new_n327_));
  INV_X1    g126(.A(G148gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .A4(KEYINPUT85), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330_));
  OAI22_X1  g129(.A1(new_n330_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G155gat), .B(G162gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n327_), .A2(new_n328_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n338_), .A2(new_n323_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n252_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(G228gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(G228gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n252_), .A2(new_n343_), .A3(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G78gat), .B(G106gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT90), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G22gat), .B(G50gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT28), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n359_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n353_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n352_), .B1(new_n252_), .B2(new_n343_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n354_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n358_), .A2(new_n362_), .B1(new_n365_), .B2(new_n356_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n356_), .A3(KEYINPUT90), .A4(new_n362_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n320_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n358_), .A2(new_n362_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n356_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n318_), .A2(new_n319_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  INV_X1    g175(.A(new_n341_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n335_), .B1(new_n325_), .B2(new_n333_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n308_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(KEYINPUT4), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n342_), .A2(KEYINPUT97), .A3(new_n381_), .A4(new_n308_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n337_), .A2(new_n341_), .A3(new_n305_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n383_), .A3(KEYINPUT4), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT96), .Z(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(new_n383_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n390_), .A2(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G85gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT0), .B(G57gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n388_), .A2(new_n398_), .A3(new_n391_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(KEYINPUT99), .A3(new_n399_), .ZN(new_n400_));
  OR3_X1    g199(.A1(new_n392_), .A2(KEYINPUT99), .A3(new_n396_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n296_), .A2(new_n375_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n373_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT32), .B(new_n280_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n280_), .A2(KEYINPUT32), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n269_), .A2(new_n406_), .A3(new_n274_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n400_), .A2(new_n401_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n397_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n392_), .A2(KEYINPUT33), .A3(new_n396_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n396_), .B1(new_n390_), .B2(new_n387_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n387_), .B2(new_n385_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n283_), .A2(new_n410_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n404_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n403_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT12), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT7), .ZN(new_n418_));
  INV_X1    g217(.A(G99gat), .ZN(new_n419_));
  INV_X1    g218(.A(G106gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n425_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n424_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n423_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G85gat), .B(G92gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT8), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n421_), .A2(new_n422_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n424_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n424_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT8), .ZN(new_n441_));
  INV_X1    g240(.A(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  OR2_X1    g242(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445_));
  NAND2_X1  g244(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n420_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT9), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G85gat), .A3(G92gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n435_), .B2(new_n450_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n433_), .B2(new_n430_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n436_), .A2(new_n443_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT66), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G78gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT11), .ZN(new_n458_));
  XOR2_X1   g257(.A(G71gat), .B(G78gat), .Z(new_n459_));
  INV_X1    g258(.A(G64gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G57gat), .ZN(new_n461_));
  INV_X1    g260(.A(G57gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G64gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n463_), .A3(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n455_), .B(new_n458_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n463_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT11), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n464_), .A3(new_n459_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n455_), .B1(new_n472_), .B2(new_n458_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n417_), .B1(new_n454_), .B2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(G230gat), .A2(G233gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n454_), .B2(new_n474_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n453_), .A2(new_n449_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT67), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n434_), .A2(KEYINPUT8), .A3(new_n435_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n441_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n436_), .A2(KEYINPUT67), .A3(new_n443_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n479_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n458_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT68), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT12), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n475_), .B(new_n477_), .C1(new_n485_), .C2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n454_), .A2(new_n474_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n454_), .A2(new_n474_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n476_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G120gat), .B(G148gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT5), .ZN(new_n496_));
  XOR2_X1   g295(.A(G176gat), .B(G204gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT13), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(KEYINPUT13), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G36gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G29gat), .ZN(new_n510_));
  INV_X1    g309(.A(G29gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G36gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n512_), .A3(KEYINPUT70), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT70), .B1(new_n510_), .B2(new_n512_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n508_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n512_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT70), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n513_), .A3(new_n507_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  INV_X1    g322(.A(G8gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n521_), .A2(new_n528_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n521_), .A2(new_n528_), .A3(KEYINPUT78), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n516_), .A2(KEYINPUT15), .A3(new_n520_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT15), .B1(new_n516_), .B2(new_n520_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n528_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(new_n534_), .A3(new_n529_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n536_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT79), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G169gat), .B(G197gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n536_), .A2(new_n540_), .A3(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n506_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n416_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G127gat), .B(G155gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT17), .Z(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n528_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n474_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n559_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT68), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n486_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n561_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n569_));
  NOR3_X1   g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n558_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n436_), .A2(KEYINPUT67), .A3(new_n443_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT67), .B1(new_n436_), .B2(new_n443_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n478_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n537_), .A2(new_n538_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n516_), .A2(new_n520_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n478_), .B(new_n579_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n436_), .A2(new_n443_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(KEYINPUT71), .A3(new_n478_), .A4(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT34), .Z(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  AND3_X1   g388(.A1(new_n578_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n575_), .A2(new_n577_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n587_), .A2(new_n588_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT71), .B1(new_n454_), .B2(new_n579_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n584_), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n597_), .A2(new_n598_), .B1(new_n485_), .B2(new_n576_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT72), .B1(new_n599_), .B2(new_n594_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n591_), .B1(new_n596_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT73), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n591_), .B(new_n609_), .C1(new_n596_), .C2(new_n600_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n610_), .A2(KEYINPUT74), .B1(new_n601_), .B2(new_n605_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n593_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n599_), .A2(KEYINPUT72), .A3(new_n594_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT74), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n591_), .A4(new_n609_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n613_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n612_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n610_), .A2(KEYINPUT74), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n606_), .A3(new_n619_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT37), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT75), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n572_), .B1(new_n622_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n553_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n402_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n523_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT38), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n552_), .A2(new_n572_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n609_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n634_), .B(new_n590_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n605_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n617_), .B2(new_n591_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n415_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n296_), .A2(new_n375_), .A3(new_n402_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n633_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n402_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT101), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n632_), .A2(new_n644_), .ZN(G1324gat));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n296_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n524_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT102), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(KEYINPUT102), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(KEYINPUT39), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n629_), .A2(new_n524_), .A3(new_n647_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n650_), .A2(KEYINPUT40), .A3(new_n652_), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n642_), .B2(new_n373_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT41), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n320_), .A2(new_n313_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n628_), .B2(new_n661_), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n366_), .A2(new_n368_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT103), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G22gat), .B1(new_n642_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n665_), .A2(G22gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n628_), .B2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n612_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n624_), .A2(new_n621_), .A3(KEYINPUT37), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n626_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n672_), .B2(new_n416_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT43), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT104), .B(new_n675_), .C1(new_n672_), .C2(new_n416_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n674_), .A2(new_n572_), .A3(new_n551_), .A4(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n571_), .B1(new_n673_), .B2(KEYINPUT43), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n551_), .A4(new_n676_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n682_), .A2(new_n511_), .A3(new_n402_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n611_), .A2(new_n571_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n553_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n630_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n683_), .A2(new_n688_), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n679_), .A2(new_n647_), .A3(new_n681_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G36gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n685_), .B(KEYINPUT105), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n296_), .B(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n509_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT45), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n687_), .A2(new_n697_), .A3(new_n509_), .A4(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n691_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n691_), .A2(new_n699_), .A3(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  OAI21_X1  g503(.A(new_n298_), .B1(new_n692_), .B2(new_n373_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n320_), .A2(G43gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n682_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g507(.A(new_n663_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G50gat), .B1(new_n682_), .B2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n665_), .A2(G50gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT107), .Z(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n692_), .B2(new_n712_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n506_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n416_), .A2(new_n549_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n627_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT108), .Z(new_n717_));
  AOI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n630_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n714_), .A2(new_n549_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n641_), .A2(new_n571_), .A3(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT109), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n462_), .B1(new_n630_), .B2(KEYINPUT110), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(KEYINPUT110), .B2(new_n462_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n721_), .B2(new_n723_), .ZN(G1332gat));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n694_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G64gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT111), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n728_), .A3(G64gat), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n727_), .A2(KEYINPUT48), .A3(new_n729_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n717_), .A2(new_n460_), .A3(new_n694_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n717_), .A2(new_n736_), .A3(new_n320_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n721_), .B2(new_n320_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n721_), .B2(new_n664_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT50), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n717_), .A2(new_n743_), .A3(new_n664_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1335gat));
  NAND4_X1  g546(.A1(new_n674_), .A2(new_n572_), .A3(new_n676_), .A4(new_n719_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n680_), .A2(new_n750_), .A3(new_n676_), .A4(new_n719_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n402_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n715_), .A2(new_n684_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n402_), .A2(G85gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(G1336gat));
  OAI21_X1  g555(.A(G92gat), .B1(new_n752_), .B2(new_n693_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n296_), .A2(G92gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n754_), .B2(new_n758_), .ZN(G1337gat));
  INV_X1    g558(.A(new_n754_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n320_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n373_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n419_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n761_), .C1(new_n762_), .C2(new_n419_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1338gat));
  NOR3_X1   g566(.A1(new_n754_), .A2(G106gat), .A3(new_n709_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G106gat), .B1(new_n748_), .B2(new_n709_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT52), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(G106gat), .C1(new_n748_), .C2(new_n709_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n768_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n768_), .B(new_n776_), .C1(new_n770_), .C2(new_n772_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  NAND3_X1  g577(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n539_), .A2(new_n535_), .A3(new_n529_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n546_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n548_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT116), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n548_), .A2(new_n781_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n499_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n490_), .B(new_n475_), .C1(new_n485_), .C2(new_n488_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n476_), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n789_));
  NAND2_X1  g588(.A1(new_n489_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n567_), .A2(new_n417_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n575_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n475_), .A4(new_n477_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n788_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n498_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n498_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(KEYINPUT118), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n786_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT58), .B(new_n786_), .C1(new_n797_), .C2(new_n800_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n622_), .A2(new_n626_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n550_), .A2(new_n499_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n796_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n500_), .A2(new_n501_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n638_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n806_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n798_), .A2(new_n799_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n795_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n810_), .B1(new_n816_), .B2(new_n807_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n817_), .C2(new_n638_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n805_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n571_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n805_), .A2(new_n819_), .A3(KEYINPUT119), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n506_), .A2(new_n549_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n672_), .A2(new_n571_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT54), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n627_), .A2(new_n827_), .A3(new_n824_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n822_), .A2(new_n823_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n296_), .A2(new_n709_), .A3(new_n320_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n402_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n826_), .A2(new_n828_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n820_), .A2(new_n572_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n831_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n550_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n820_), .A2(new_n821_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n572_), .A3(new_n823_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n832_), .B1(new_n842_), .B2(new_n834_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n550_), .A2(G113gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n844_), .B2(new_n845_), .ZN(G1340gat));
  OAI211_X1 g645(.A(new_n506_), .B(new_n838_), .C1(new_n843_), .C2(new_n837_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT120), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n833_), .A2(new_n849_), .A3(new_n506_), .A4(new_n838_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(G120gat), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n714_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n843_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n844_), .B2(new_n572_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT121), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n856_), .C1(new_n844_), .C2(new_n572_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n839_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n571_), .A2(G127gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT122), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n858_), .A2(new_n860_), .B1(new_n861_), .B2(new_n863_), .ZN(G1342gat));
  OAI21_X1  g663(.A(G134gat), .B1(new_n839_), .B2(new_n672_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n611_), .A2(G134gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n844_), .B2(new_n866_), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n842_), .A2(new_n834_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n694_), .A2(new_n402_), .A3(new_n374_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n550_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n327_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n714_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n328_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n870_), .A2(new_n572_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n870_), .B2(new_n672_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n611_), .A2(G162gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n870_), .B2(new_n879_), .ZN(G1347gat));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n664_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n693_), .A2(new_n630_), .A3(new_n373_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n550_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n881_), .B1(new_n885_), .B2(new_n216_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n203_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT62), .B(G169gat), .C1(new_n884_), .C2(new_n550_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(G1348gat));
  OAI21_X1  g688(.A(new_n204_), .B1(new_n884_), .B2(new_n714_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n892_), .B(new_n204_), .C1(new_n884_), .C2(new_n714_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n829_), .A2(new_n663_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n883_), .A2(G176gat), .A3(new_n506_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n891_), .A2(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n883_), .A2(new_n571_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n882_), .A2(new_n264_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n898_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n208_), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n884_), .B2(new_n672_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n611_), .A2(new_n263_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n884_), .B2(new_n903_), .ZN(G1351gat));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT124), .B1(new_n630_), .B2(new_n374_), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n630_), .A2(KEYINPUT124), .A3(new_n374_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n694_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n905_), .B1(new_n829_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n908_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n868_), .A2(KEYINPUT125), .A3(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n550_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT126), .B(G197gat), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n912_), .B(new_n914_), .ZN(G1352gat));
  AOI21_X1  g714(.A(new_n714_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n238_), .ZN(G1353gat));
  NAND2_X1  g716(.A1(new_n909_), .A2(new_n911_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n572_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n918_), .A2(new_n922_), .A3(new_n919_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1354gat));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n918_), .A2(new_n927_), .A3(new_n638_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n672_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n927_), .ZN(G1355gat));
endmodule


