//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT74), .ZN(new_n203_));
  XOR2_X1   g002(.A(G43gat), .B(G50gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n211_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT8), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n210_), .B1(new_n209_), .B2(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n208_), .A2(KEYINPUT65), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(new_n208_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n220_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT66), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n220_), .B(new_n226_), .C1(new_n223_), .C2(new_n222_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n217_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT10), .B(G99gat), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n234_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n228_), .B(new_n229_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n219_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n229_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT70), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n207_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT76), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n218_), .B(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n245_), .B2(new_n240_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(new_n247_), .A3(new_n219_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n205_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(KEYINPUT76), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n243_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G232gat), .A2(G233gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT34), .Z(new_n254_));
  XNOR2_X1  g053(.A(G190gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G134gat), .B(G162gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n252_), .A2(new_n254_), .B1(KEYINPUT36), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n254_), .B(KEYINPUT73), .Z(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT35), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n252_), .B2(KEYINPUT77), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n251_), .A2(new_n250_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n243_), .A4(new_n260_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n257_), .A2(KEYINPUT36), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n258_), .A2(new_n262_), .A3(new_n269_), .A4(new_n265_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT37), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(KEYINPUT37), .A3(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G127gat), .B(G155gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT16), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G183gat), .B(G211gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT17), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n280_), .A2(KEYINPUT80), .A3(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G1gat), .B(G8gat), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT78), .B(G15gat), .ZN(new_n285_));
  INV_X1    g084(.A(G22gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n288_));
  INV_X1    g087(.A(G1gat), .ZN(new_n289_));
  INV_X1    g088(.A(G8gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT14), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n287_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n284_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n283_), .A3(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G71gat), .B(G78gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n302_), .A2(new_n304_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n300_), .B(new_n309_), .ZN(new_n310_));
  AOI211_X1 g109(.A(new_n282_), .B(new_n310_), .C1(new_n281_), .C2(new_n280_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n282_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT81), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n276_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT94), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT19), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT21), .ZN(new_n321_));
  INV_X1    g120(.A(G218gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G211gat), .ZN(new_n323_));
  INV_X1    g122(.A(G211gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G218gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G204gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT91), .B1(new_n327_), .B2(G197gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(G204gat), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n330_), .B2(G204gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n326_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT92), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n329_), .B1(new_n330_), .B2(G204gat), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n327_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n334_), .B(new_n335_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n326_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n330_), .B2(G204gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n327_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n330_), .A2(G204gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT21), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n323_), .A2(new_n325_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n350_), .B(new_n351_), .C1(new_n341_), .C2(KEYINPUT21), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT25), .B(G183gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT24), .ZN(new_n361_));
  INV_X1    g160(.A(G169gat), .ZN(new_n362_));
  INV_X1    g161(.A(G176gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT24), .A3(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n355_), .A2(new_n360_), .A3(new_n364_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(G169gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G169gat), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n363_), .B(new_n371_), .C1(new_n372_), .C2(new_n369_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n358_), .B(new_n359_), .C1(G183gat), .C2(G190gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n366_), .A3(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n344_), .A2(new_n352_), .A3(new_n368_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n363_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n374_), .A3(new_n366_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n368_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n344_), .B2(new_n352_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT20), .B(new_n376_), .C1(new_n380_), .C2(KEYINPUT93), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n341_), .A2(new_n342_), .A3(new_n326_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n342_), .B1(new_n341_), .B2(new_n326_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n352_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n368_), .A2(new_n378_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n318_), .B(new_n320_), .C1(new_n381_), .C2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n320_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n375_), .A2(new_n368_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT93), .B1(new_n384_), .B2(new_n385_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n386_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n388_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n384_), .A2(new_n389_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n344_), .A2(new_n352_), .A3(new_n379_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT20), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT94), .B1(new_n397_), .B2(new_n320_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n387_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n387_), .B(new_n406_), .C1(new_n394_), .C2(new_n398_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n317_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n399_), .A2(new_n404_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n392_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n397_), .A2(new_n320_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n413_), .A2(KEYINPUT101), .A3(new_n406_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT101), .B1(new_n413_), .B2(new_n406_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT27), .B(new_n410_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(KEYINPUT1), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(KEYINPUT1), .B2(new_n419_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G141gat), .A2(G148gat), .ZN(new_n422_));
  INV_X1    g221(.A(G141gat), .ZN(new_n423_));
  INV_X1    g222(.A(G148gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n422_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT2), .ZN(new_n428_));
  OR3_X1    g227(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT87), .B(KEYINPUT2), .Z(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT88), .A3(new_n422_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n427_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n431_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n418_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n419_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n426_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  OR3_X1    g239(.A1(new_n440_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT28), .B1(new_n440_), .B2(KEYINPUT29), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(KEYINPUT29), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n384_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n384_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G228gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G78gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(new_n232_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G22gat), .B(G50gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n445_), .A2(new_n447_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n417_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G134gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G127gat), .ZN(new_n460_));
  INV_X1    g259(.A(G127gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G134gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n462_), .A3(KEYINPUT86), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G113gat), .B(G120gat), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n467_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n470_), .B(new_n426_), .C1(new_n437_), .C2(new_n439_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n468_), .A2(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n440_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT97), .A4(new_n474_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT4), .ZN(new_n480_));
  INV_X1    g279(.A(new_n474_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n440_), .A2(new_n472_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G85gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT100), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n477_), .A3(new_n489_), .A4(new_n478_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n485_), .A2(KEYINPUT100), .A3(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G43gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT30), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(new_n389_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT85), .B(G15gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n472_), .B(KEYINPUT31), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G227gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n506_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n497_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n458_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n456_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n512_), .A2(new_n409_), .A3(new_n416_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT98), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n410_), .A2(new_n515_), .A3(new_n407_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n479_), .A2(new_n517_), .A3(new_n489_), .A4(new_n484_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n493_), .A2(KEYINPUT33), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n480_), .A2(new_n474_), .A3(new_n483_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n471_), .A2(new_n473_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n489_), .B1(new_n521_), .B2(new_n481_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n518_), .A2(new_n519_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n515_), .B1(new_n410_), .B2(new_n407_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n514_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT96), .B1(new_n405_), .B2(new_n408_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n527_), .A2(KEYINPUT98), .A3(new_n516_), .A4(new_n523_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n411_), .A2(new_n412_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT99), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n399_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n399_), .B2(KEYINPUT99), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n494_), .B(new_n495_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n513_), .B1(new_n535_), .B2(new_n456_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n509_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n511_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n295_), .A2(new_n297_), .A3(new_n205_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n205_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n541_));
  OAI211_X1 g340(.A(G229gat), .B(G233gat), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n207_), .A2(new_n298_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT82), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G113gat), .B(G141gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT83), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G169gat), .B(G197gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n546_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n538_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n309_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n249_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT68), .A4(new_n309_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n246_), .A2(new_n248_), .A3(new_n309_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT68), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n559_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT12), .B(new_n309_), .C1(new_n238_), .C2(new_n241_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n561_), .A3(new_n570_), .A4(new_n558_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(KEYINPUT69), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(KEYINPUT69), .B2(new_n567_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT71), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n316_), .A2(new_n557_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n289_), .A3(new_n497_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n556_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n313_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n538_), .A2(new_n271_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n496_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n587_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n417_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(G8gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n585_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G8gat), .B1(new_n594_), .B2(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT102), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n602_), .B2(KEYINPUT39), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n601_), .A2(KEYINPUT102), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(KEYINPUT39), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n604_), .B(KEYINPUT40), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n605_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n603_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(G1325gat));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n593_), .B2(new_n537_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n585_), .A2(new_n612_), .A3(new_n537_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  AOI21_X1  g415(.A(new_n286_), .B1(new_n593_), .B2(new_n457_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT42), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n585_), .A2(new_n286_), .A3(new_n457_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1327gat));
  NOR2_X1   g419(.A1(new_n314_), .A2(new_n271_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n557_), .A2(new_n584_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(G29gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n497_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n535_), .A2(new_n456_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n513_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n537_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n511_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n625_), .B(new_n275_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT103), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n538_), .A2(new_n632_), .A3(new_n625_), .A4(new_n275_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n538_), .A2(new_n275_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT43), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n589_), .A2(new_n314_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n637_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n497_), .A3(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n642_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT104), .B1(new_n642_), .B2(G29gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n624_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT105), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(new_n624_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n622_), .A2(new_n650_), .A3(new_n417_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT45), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n640_), .A2(new_n417_), .A3(new_n641_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n653_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT106), .B1(new_n653_), .B2(G36gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n652_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT46), .B(new_n652_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  AOI21_X1  g459(.A(G43gat), .B1(new_n622_), .B2(new_n537_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n640_), .A2(new_n641_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n537_), .A2(G43gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g464(.A(G50gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n622_), .A2(new_n666_), .A3(new_n457_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(KEYINPUT107), .A3(new_n457_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT107), .B1(new_n662_), .B2(new_n457_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(G1331gat));
  NOR2_X1   g470(.A1(new_n584_), .A2(new_n556_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n538_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n316_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n496_), .B1(new_n674_), .B2(KEYINPUT108), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(KEYINPUT108), .B2(new_n674_), .ZN(new_n676_));
  INV_X1    g475(.A(G57gat), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n592_), .A2(new_n314_), .A3(new_n672_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n496_), .A2(new_n677_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n676_), .A2(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(G1332gat));
  INV_X1    g479(.A(G64gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n678_), .B2(new_n417_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT48), .Z(new_n683_));
  INV_X1    g482(.A(new_n674_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n681_), .A3(new_n417_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1333gat));
  INV_X1    g487(.A(G71gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n678_), .B2(new_n537_), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n537_), .A2(new_n689_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n674_), .B2(new_n693_), .ZN(G1334gat));
  AOI21_X1  g493(.A(new_n449_), .B1(new_n678_), .B2(new_n457_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT50), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n449_), .A3(new_n457_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1335gat));
  AND2_X1   g497(.A1(new_n673_), .A2(new_n621_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G85gat), .B1(new_n699_), .B2(new_n497_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT111), .ZN(new_n701_));
  INV_X1    g500(.A(new_n314_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n636_), .A2(new_n702_), .A3(new_n672_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n497_), .A2(G85gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(G1336gat));
  INV_X1    g504(.A(G92gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n706_), .A3(new_n417_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n703_), .A2(new_n417_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(new_n706_), .ZN(G1337gat));
  NAND2_X1  g508(.A1(new_n703_), .A2(new_n537_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G99gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n699_), .A2(new_n537_), .A3(new_n231_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT113), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n714_), .B(new_n716_), .Z(G1338gat));
  NAND3_X1  g516(.A1(new_n699_), .A2(new_n232_), .A3(new_n457_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n636_), .A2(new_n457_), .A3(new_n702_), .A4(new_n672_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .A4(G106gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n232_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n720_), .A2(new_n723_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g525(.A(KEYINPUT122), .ZN(new_n727_));
  INV_X1    g526(.A(G113gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n458_), .A2(new_n497_), .A3(new_n537_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n559_), .A2(KEYINPUT116), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n569_), .A2(new_n561_), .A3(new_n570_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n559_), .A2(KEYINPUT55), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n731_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n569_), .A2(new_n561_), .A3(new_n570_), .A4(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n571_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n734_), .A2(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n571_), .A2(KEYINPUT115), .A3(new_n737_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n578_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(KEYINPUT56), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n555_), .B1(new_n573_), .B2(new_n578_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT118), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n734_), .A2(new_n736_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n738_), .A2(new_n739_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n741_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n578_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n743_), .B2(KEYINPUT56), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n755_), .A2(new_n745_), .A3(new_n756_), .A4(new_n747_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT119), .ZN(new_n758_));
  INV_X1    g557(.A(new_n545_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n541_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n539_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n761_), .B2(new_n551_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n545_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(KEYINPUT119), .A3(new_n550_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n543_), .A2(new_n539_), .A3(new_n759_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n552_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(KEYINPUT120), .A3(new_n552_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n580_), .A2(new_n771_), .A3(new_n581_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n749_), .A2(new_n757_), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT57), .A3(new_n271_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT121), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n774_), .A2(new_n777_), .A3(KEYINPUT57), .A4(new_n271_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n769_), .A2(new_n770_), .B1(new_n573_), .B2(new_n578_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .A4(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n275_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n774_), .A2(new_n271_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n313_), .B1(new_n779_), .B2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n276_), .A2(new_n314_), .A3(new_n555_), .A4(new_n584_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT54), .Z(new_n794_));
  OAI21_X1  g593(.A(new_n730_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n793_), .B(KEYINPUT54), .ZN(new_n796_));
  INV_X1    g595(.A(new_n271_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n755_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n772_), .B1(new_n798_), .B2(KEYINPUT118), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(new_n757_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n787_), .B1(new_n800_), .B2(KEYINPUT57), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n796_), .B1(new_n802_), .B2(new_n314_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n729_), .A2(KEYINPUT59), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n795_), .A2(KEYINPUT59), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n728_), .B1(new_n805_), .B2(new_n556_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n795_), .A2(G113gat), .A3(new_n555_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n727_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n804_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n779_), .A2(new_n791_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n590_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n729_), .B1(new_n811_), .B2(new_n796_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n809_), .B(new_n556_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G113gat), .ZN(new_n815_));
  INV_X1    g614(.A(new_n807_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT122), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n808_), .A2(new_n817_), .ZN(G1340gat));
  INV_X1    g617(.A(new_n805_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G120gat), .B1(new_n819_), .B2(new_n584_), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n584_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(KEYINPUT60), .B2(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n820_), .B1(new_n795_), .B2(new_n823_), .ZN(G1341gat));
  OAI21_X1  g623(.A(G127gat), .B1(new_n819_), .B2(new_n590_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n812_), .A2(new_n461_), .A3(new_n314_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1342gat));
  OAI21_X1  g626(.A(G134gat), .B1(new_n819_), .B2(new_n276_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n812_), .A2(new_n459_), .A3(new_n797_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n811_), .A2(new_n796_), .ZN(new_n831_));
  NOR4_X1   g630(.A1(new_n417_), .A2(new_n496_), .A3(new_n456_), .A4(new_n537_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT123), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n555_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(new_n423_), .ZN(G1344gat));
  NOR2_X1   g635(.A1(new_n834_), .A2(new_n584_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(new_n424_), .ZN(G1345gat));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n702_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT61), .B(G155gat), .Z(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  INV_X1    g640(.A(new_n834_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G162gat), .B1(new_n842_), .B2(new_n797_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n275_), .A2(G162gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT124), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n842_), .B2(new_n845_), .ZN(G1347gat));
  INV_X1    g645(.A(KEYINPUT126), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n510_), .A2(new_n417_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT125), .Z(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n457_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n803_), .A2(new_n556_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n803_), .A2(new_n372_), .A3(new_n556_), .A4(new_n850_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT62), .B1(new_n851_), .B2(G169gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n847_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n855_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(KEYINPUT126), .A3(new_n853_), .A4(new_n852_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1348gat));
  NAND2_X1  g658(.A1(new_n803_), .A2(new_n850_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n584_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G176gat), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n457_), .B1(new_n811_), .B2(new_n796_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n849_), .A2(new_n584_), .A3(new_n363_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1349gat));
  NOR3_X1   g665(.A1(new_n860_), .A2(new_n353_), .A3(new_n590_), .ZN(new_n867_));
  INV_X1    g666(.A(G183gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n849_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n314_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n868_), .B2(new_n870_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n860_), .B2(new_n276_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n797_), .A2(new_n354_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n860_), .B2(new_n873_), .ZN(G1351gat));
  AND3_X1   g673(.A1(new_n417_), .A2(new_n512_), .A3(new_n509_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n831_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n555_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n330_), .ZN(G1352gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n584_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n327_), .ZN(G1353gat));
  NOR2_X1   g679(.A1(new_n876_), .A2(new_n590_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n881_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT63), .B(G211gat), .Z(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(new_n883_), .ZN(G1354gat));
  NOR3_X1   g683(.A1(new_n876_), .A2(new_n322_), .A3(new_n276_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n876_), .A2(new_n271_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT127), .ZN(new_n887_));
  AOI21_X1  g686(.A(G218gat), .B1(new_n886_), .B2(KEYINPUT127), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n885_), .B1(new_n887_), .B2(new_n888_), .ZN(G1355gat));
endmodule


