//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_;
  INV_X1    g000(.A(G230gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n206_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n211_), .A2(KEYINPUT65), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(G99gat), .A4(G106gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT64), .B(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT65), .B1(new_n211_), .B2(new_n213_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n214_), .A2(new_n224_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n230_), .A2(new_n231_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n220_), .B(new_n223_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n209_), .A2(new_n210_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n229_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n247_), .B(new_n229_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n205_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT68), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n240_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n254_), .A3(KEYINPUT12), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n240_), .B(new_n248_), .C1(new_n253_), .C2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n205_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT70), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n261_), .A3(new_n205_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n258_), .A2(new_n263_), .A3(KEYINPUT71), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT71), .B1(new_n258_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n252_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G120gat), .B(G148gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(G176gat), .B(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n252_), .B(new_n273_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(KEYINPUT73), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n266_), .A2(new_n276_), .A3(new_n271_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT13), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT75), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n285_));
  XOR2_X1   g084(.A(G29gat), .B(G36gat), .Z(new_n286_));
  INV_X1    g085(.A(G43gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G29gat), .B(G36gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G43gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(G50gat), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(G50gat), .B1(new_n288_), .B2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n285_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(KEYINPUT80), .A3(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  INV_X1    g097(.A(G1gat), .ZN(new_n299_));
  INV_X1    g098(.A(G8gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT14), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G8gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT81), .B1(new_n297_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT81), .ZN(new_n307_));
  AOI211_X1 g106(.A(new_n307_), .B(new_n304_), .C1(new_n294_), .C2(new_n296_), .ZN(new_n308_));
  OAI22_X1  g107(.A1(new_n306_), .A2(new_n308_), .B1(new_n305_), .B2(new_n297_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n292_), .A2(new_n293_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(KEYINPUT15), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(KEYINPUT15), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n304_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(new_n310_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G141gat), .ZN(new_n318_));
  INV_X1    g117(.A(G169gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(G197gat), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT82), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n312_), .A2(new_n325_), .A3(new_n317_), .A4(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n312_), .A2(new_n317_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n321_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G183gat), .ZN(new_n332_));
  INV_X1    g131(.A(G190gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT23), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  MUX2_X1   g136(.A(new_n337_), .B(new_n336_), .S(KEYINPUT85), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT25), .B(G183gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT84), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G176gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n319_), .B2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(KEYINPUT24), .ZN(new_n347_));
  INV_X1    g146(.A(new_n344_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT24), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n338_), .B(new_n341_), .C1(new_n347_), .C2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n337_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT98), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n319_), .A2(new_n345_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G169gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n345_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G197gat), .B(G204gat), .Z(new_n358_));
  AND2_X1   g157(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n358_), .B2(KEYINPUT21), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n361_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT99), .B1(new_n357_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT97), .Z(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT19), .Z(new_n368_));
  OAI21_X1  g167(.A(new_n338_), .B1(G183gat), .B2(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n355_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n347_), .A2(new_n349_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n333_), .A2(KEYINPUT26), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n340_), .B1(KEYINPUT83), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n339_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n337_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n370_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n368_), .B1(new_n377_), .B2(new_n364_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n364_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT99), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n350_), .A2(new_n379_), .A3(new_n356_), .A4(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n365_), .A2(new_n378_), .A3(KEYINPUT20), .A4(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT20), .B1(new_n377_), .B2(new_n364_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n368_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n382_), .A2(new_n385_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT101), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n386_), .A2(KEYINPUT101), .A3(new_n391_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT91), .ZN(new_n399_));
  NOR3_X1   g198(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(KEYINPUT90), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(KEYINPUT90), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT2), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(KEYINPUT92), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT92), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(KEYINPUT1), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n406_), .B(KEYINPUT88), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT1), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n418_), .A3(new_n409_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G141gat), .B(G148gat), .Z(new_n420_));
  AND3_X1   g219(.A1(new_n419_), .A2(KEYINPUT89), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT89), .B1(new_n419_), .B2(new_n420_), .ZN(new_n422_));
  OAI22_X1  g221(.A1(new_n412_), .A2(new_n414_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G127gat), .B(G134gat), .ZN(new_n424_));
  INV_X1    g223(.A(G113gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G120gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n411_), .B(KEYINPUT92), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n419_), .A2(new_n420_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n419_), .A2(KEYINPUT89), .A3(new_n420_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n436_), .A3(new_n428_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n437_), .A3(KEYINPUT4), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT102), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT102), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n430_), .A2(new_n437_), .A3(new_n440_), .A4(KEYINPUT4), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(new_n430_), .B2(KEYINPUT4), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n423_), .A2(KEYINPUT103), .A3(new_n444_), .A4(new_n429_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n439_), .A2(new_n441_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT0), .B(G57gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G85gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(G1gat), .B(G29gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n430_), .A2(new_n437_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n447_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n396_), .A2(new_n397_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n447_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n459_), .B1(new_n446_), .B2(new_n454_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n460_), .B2(new_n452_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n439_), .A2(new_n441_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n443_), .A2(new_n445_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n454_), .A3(new_n463_), .ZN(new_n464_));
  AND4_X1   g263(.A1(new_n457_), .A2(new_n464_), .A3(new_n458_), .A4(new_n452_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n456_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT104), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n468_));
  INV_X1    g267(.A(new_n368_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n364_), .B(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n350_), .A2(new_n356_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n474_), .A2(KEYINPUT105), .B1(new_n377_), .B2(new_n364_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n364_), .B(KEYINPUT95), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT20), .B1(new_n476_), .B2(new_n357_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT105), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n469_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n383_), .A2(new_n368_), .A3(new_n384_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n468_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n460_), .A2(new_n452_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n460_), .A2(new_n452_), .ZN(new_n484_));
  OAI221_X1 g283(.A(new_n482_), .B1(new_n386_), .B2(new_n468_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT104), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n456_), .C1(new_n461_), .C2(new_n465_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n467_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n428_), .B(KEYINPUT31), .Z(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT87), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(new_n377_), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G43gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G15gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n493_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G71gat), .B(G99gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n491_), .B(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n500_));
  OR3_X1    g299(.A1(new_n423_), .A2(KEYINPUT29), .A3(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n423_), .B2(KEYINPUT29), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G22gat), .B(G50gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT96), .ZN(new_n506_));
  NAND2_X1  g305(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(G228gat), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n423_), .A2(KEYINPUT29), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n511_), .B2(new_n476_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n379_), .B1(new_n423_), .B2(KEYINPUT29), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G78gat), .B(G106gat), .Z(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n515_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n505_), .B1(new_n520_), .B2(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT96), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n488_), .A2(new_n499_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n499_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n519_), .A2(new_n499_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n483_), .A2(new_n484_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT27), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n396_), .A2(new_n530_), .A3(new_n397_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT107), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n394_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n480_), .A2(new_n481_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n393_), .A2(KEYINPUT106), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n393_), .A2(KEYINPUT106), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n533_), .A2(new_n534_), .B1(new_n540_), .B2(KEYINPUT27), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n528_), .A2(new_n529_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n331_), .B1(new_n524_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n284_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n529_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n313_), .B(KEYINPUT15), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(new_n240_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT34), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT77), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n313_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n240_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n551_), .A2(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT76), .B(G134gat), .ZN(new_n559_));
  INV_X1    g358(.A(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT36), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n548_), .A2(new_n555_), .B1(new_n552_), .B2(new_n551_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n558_), .B2(new_n565_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n546_), .B(KEYINPUT37), .C1(new_n567_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n546_), .A2(KEYINPUT37), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n546_), .A2(KEYINPUT37), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n571_), .A2(new_n566_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n304_), .B(KEYINPUT79), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(new_n248_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n248_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT16), .B(G183gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT69), .A3(KEYINPUT17), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n586_), .A2(KEYINPUT17), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n579_), .A2(new_n580_), .B1(new_n589_), .B2(new_n587_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n575_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n544_), .A2(new_n299_), .A3(new_n545_), .A4(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n283_), .A2(new_n543_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n567_), .A2(new_n569_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n591_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n545_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G1gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n593_), .A2(new_n594_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(G1324gat));
  NOR2_X1   g402(.A1(new_n541_), .A2(G8gat), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n284_), .A2(new_n543_), .A3(new_n592_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n541_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n283_), .A2(new_n543_), .A3(new_n599_), .A4(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n607_), .A2(new_n608_), .A3(G8gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n607_), .B2(G8gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n605_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT109), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT109), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n605_), .B(new_n613_), .C1(new_n610_), .C2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT40), .ZN(G1325gat));
  NAND3_X1  g415(.A1(new_n596_), .A2(new_n599_), .A3(new_n525_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(G15gat), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT41), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G15gat), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n544_), .A2(new_n621_), .A3(new_n525_), .A4(new_n592_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT110), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n523_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n544_), .A2(new_n626_), .A3(new_n627_), .A4(new_n592_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n596_), .A2(new_n599_), .A3(new_n627_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G22gat), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(KEYINPUT42), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(KEYINPUT42), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT111), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1327gat));
  NAND2_X1  g434(.A1(new_n524_), .A2(new_n542_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n575_), .B(KEYINPUT112), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT43), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n575_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n524_), .B2(new_n542_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n331_), .B1(new_n639_), .B2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n591_), .A4(new_n283_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n640_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n591_), .B(new_n330_), .C1(new_n647_), .C2(new_n642_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n283_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n650_), .ZN(new_n651_));
  OR3_X1    g450(.A1(new_n651_), .A2(KEYINPUT113), .A3(new_n529_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT113), .B1(new_n651_), .B2(new_n529_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(G29gat), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n591_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n597_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n283_), .A2(new_n543_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n529_), .A2(G29gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT114), .Z(new_n660_));
  OAI21_X1  g459(.A(new_n654_), .B1(new_n658_), .B2(new_n660_), .ZN(G1328gat));
  OAI21_X1  g460(.A(G36gat), .B1(new_n651_), .B2(new_n541_), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n663_), .A3(new_n606_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT45), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n662_), .A2(new_n665_), .A3(KEYINPUT46), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1329gat));
  INV_X1    g469(.A(KEYINPUT47), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n499_), .A2(new_n287_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n645_), .A2(new_n650_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT115), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n287_), .B1(new_n658_), .B2(new_n499_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n671_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n673_), .A2(new_n675_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT115), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(KEYINPUT47), .A3(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1330gat));
  OAI21_X1  g482(.A(G50gat), .B1(new_n651_), .B2(new_n523_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n658_), .A2(G50gat), .A3(new_n523_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1331gat));
  AOI21_X1  g485(.A(new_n330_), .B1(new_n524_), .B2(new_n542_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT116), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(new_n649_), .A3(new_n592_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G57gat), .B1(new_n689_), .B2(new_n545_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT75), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n283_), .B(new_n691_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(new_n599_), .A3(new_n687_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n545_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n690_), .B1(new_n694_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n693_), .B2(new_n606_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT48), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n689_), .A2(new_n696_), .A3(new_n606_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n693_), .B2(new_n525_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT49), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n689_), .A2(new_n701_), .A3(new_n525_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1334gat));
  INV_X1    g504(.A(G78gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n693_), .B2(new_n627_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT50), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n689_), .A2(new_n706_), .A3(new_n627_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1335gat));
  AND3_X1   g509(.A1(new_n692_), .A2(new_n656_), .A3(new_n688_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n545_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n283_), .B1(new_n639_), .B2(new_n643_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n591_), .A3(new_n331_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n714_), .A2(new_n207_), .A3(new_n529_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1336gat));
  AOI21_X1  g515(.A(G92gat), .B1(new_n711_), .B2(new_n606_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n714_), .A2(new_n208_), .A3(new_n541_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1337gat));
  INV_X1    g518(.A(KEYINPUT117), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(KEYINPUT51), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n711_), .A2(new_n225_), .A3(new_n525_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G99gat), .B1(new_n714_), .B2(new_n499_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n720_), .A2(KEYINPUT51), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n226_), .A3(new_n627_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n713_), .A2(new_n591_), .A3(new_n331_), .A4(new_n627_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(G106gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n728_), .B2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n727_), .B(new_n735_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  INV_X1    g536(.A(KEYINPUT122), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n591_), .A2(new_n330_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT118), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n575_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT118), .B1(new_n591_), .B2(new_n330_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n275_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n741_), .B(new_n742_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n258_), .A2(new_n263_), .A3(KEYINPUT55), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n258_), .A2(new_n250_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n204_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n750_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n271_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n756_), .A3(new_n271_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n755_), .A2(new_n330_), .A3(new_n274_), .A4(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n316_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT119), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT119), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n316_), .B(new_n761_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n311_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n309_), .A2(new_n310_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n765_), .A2(new_n321_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n275_), .A2(new_n766_), .A3(new_n277_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n275_), .A2(new_n766_), .A3(KEYINPUT120), .A4(new_n277_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n758_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT121), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n597_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n755_), .A2(new_n274_), .A3(new_n757_), .A4(new_n766_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n779_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n575_), .A3(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n771_), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n597_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n774_), .A2(new_n777_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n747_), .B1(new_n784_), .B2(new_n591_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n606_), .A2(new_n529_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n526_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT59), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n738_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT122), .B(KEYINPUT59), .C1(new_n785_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n747_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n784_), .A2(KEYINPUT123), .A3(new_n591_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT123), .B1(new_n784_), .B2(new_n591_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n788_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n790_), .A3(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n793_), .A2(G113gat), .A3(new_n330_), .A4(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n784_), .A2(new_n591_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n794_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n798_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n425_), .B1(new_n803_), .B2(new_n331_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1340gat));
  AOI21_X1  g604(.A(KEYINPUT122), .B1(new_n803_), .B2(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(new_n792_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n799_), .B(new_n692_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT124), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n793_), .A2(KEYINPUT124), .A3(new_n692_), .A4(new_n799_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(G120gat), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n427_), .B1(new_n283_), .B2(KEYINPUT60), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n789_), .B(new_n813_), .C1(KEYINPUT60), .C2(new_n427_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1341gat));
  AOI21_X1  g614(.A(G127gat), .B1(new_n789_), .B2(new_n655_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n793_), .A2(new_n655_), .A3(new_n799_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g617(.A(G134gat), .B1(new_n789_), .B2(new_n598_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n793_), .A2(new_n575_), .A3(new_n799_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g620(.A1(new_n785_), .A2(new_n527_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n786_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT125), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(KEYINPUT125), .A3(new_n786_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n330_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n692_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n655_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT61), .B(G155gat), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1346gat));
  AOI21_X1  g633(.A(G162gat), .B1(new_n827_), .B2(new_n598_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n560_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n637_), .B2(new_n836_), .ZN(G1347gat));
  NOR2_X1   g636(.A1(new_n541_), .A2(new_n545_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n525_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n797_), .A2(new_n330_), .A3(new_n523_), .A4(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G169gat), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n797_), .A2(new_n523_), .A3(new_n840_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n330_), .A3(new_n354_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n841_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(G1348gat));
  AOI21_X1  g647(.A(G176gat), .B1(new_n845_), .B2(new_n649_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n802_), .A2(new_n523_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n284_), .A2(new_n345_), .A3(new_n839_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(G1349gat));
  NOR2_X1   g652(.A1(new_n591_), .A2(new_n340_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n655_), .A3(new_n840_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n845_), .A2(new_n854_), .B1(new_n855_), .B2(new_n332_), .ZN(G1350gat));
  NAND3_X1  g655(.A1(new_n845_), .A2(new_n598_), .A3(new_n339_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n845_), .A2(new_n575_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n333_), .ZN(G1351gat));
  NAND2_X1  g658(.A1(new_n822_), .A2(new_n838_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n330_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g662(.A(G204gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT126), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT126), .B(G204gat), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n860_), .A2(new_n284_), .ZN(new_n867_));
  MUX2_X1   g666(.A(new_n865_), .B(new_n866_), .S(new_n867_), .Z(G1353gat));
  NAND2_X1  g667(.A1(new_n861_), .A2(new_n655_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  AND2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n869_), .B2(new_n870_), .ZN(G1354gat));
  NOR2_X1   g672(.A1(new_n860_), .A2(new_n597_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n861_), .A2(new_n575_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT127), .B(G218gat), .ZN(new_n876_));
  MUX2_X1   g675(.A(new_n874_), .B(new_n875_), .S(new_n876_), .Z(G1355gat));
endmodule


