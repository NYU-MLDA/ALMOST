//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT6), .B1(new_n206_), .B2(new_n205_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n204_), .A2(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G85gat), .Z(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(G92gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(KEYINPUT65), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n210_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G85gat), .B(G92gat), .Z(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT8), .B1(new_n220_), .B2(KEYINPUT67), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT66), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n207_), .A2(new_n209_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n223_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n219_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n207_), .A2(new_n209_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n226_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n224_), .B(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n220_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n221_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT68), .B1(new_n230_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT64), .B(G85gat), .ZN(new_n239_));
  INV_X1    g038(.A(G92gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n211_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n217_), .A3(new_n216_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n236_), .A2(new_n221_), .B1(new_n242_), .B2(new_n210_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n229_), .A2(new_n222_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G64gat), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n249_));
  XOR2_X1   g048(.A(G71gat), .B(G78gat), .Z(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n238_), .A2(new_n246_), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT69), .ZN(new_n255_));
  INV_X1    g054(.A(new_n253_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n230_), .A2(new_n237_), .A3(KEYINPUT68), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(KEYINPUT69), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n255_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n261_), .A2(KEYINPUT70), .A3(new_n263_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269_));
  OAI211_X1 g068(.A(KEYINPUT12), .B(new_n256_), .C1(new_n230_), .C2(new_n237_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n253_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n254_), .B(new_n270_), .C1(new_n271_), .C2(KEYINPUT12), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n272_), .B2(new_n263_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n254_), .A2(new_n270_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n259_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n274_), .A2(new_n276_), .A3(KEYINPUT71), .A4(new_n262_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n268_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n268_), .B2(new_n278_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n203_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT13), .A3(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n230_), .A2(new_n237_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G29gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G43gat), .B(G50gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n294_), .B(KEYINPUT15), .Z(new_n295_));
  NOR2_X1   g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n238_), .A2(new_n246_), .A3(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT34), .Z(new_n302_));
  XOR2_X1   g101(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n302_), .A2(new_n303_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n296_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n300_), .A2(new_n304_), .B1(new_n299_), .B2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G190gat), .B(G218gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(G134gat), .B(G162gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT36), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT75), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n311_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT74), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n307_), .A2(new_n312_), .ZN(new_n318_));
  OAI211_X1 g117(.A(KEYINPUT37), .B(new_n313_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n307_), .A2(new_n312_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT37), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n320_), .B(new_n316_), .C1(KEYINPUT75), .C2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G15gat), .B(G22gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(G1gat), .A2(G8gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(KEYINPUT14), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT76), .ZN(new_n328_));
  XOR2_X1   g127(.A(G1gat), .B(G8gat), .Z(new_n329_));
  OR2_X1    g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n329_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G231gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n253_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n332_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n336_));
  XOR2_X1   g135(.A(G127gat), .B(G155gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT16), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G183gat), .B(G211gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n335_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(KEYINPUT17), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n290_), .A2(new_n324_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n347_), .B(new_n348_), .C1(G183gat), .C2(G190gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G169gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G190gat), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT25), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT79), .B(KEYINPUT25), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT80), .B1(new_n360_), .B2(new_n354_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(KEYINPUT25), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT79), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n362_), .B(G183gat), .C1(new_n364_), .C2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n359_), .B1(new_n361_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369_));
  INV_X1    g168(.A(G169gat), .ZN(new_n370_));
  INV_X1    g169(.A(G176gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n347_), .A2(new_n348_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n373_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n352_), .B1(new_n368_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(G15gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT30), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n381_), .B(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G127gat), .B(G134gat), .Z(new_n387_));
  XOR2_X1   g186(.A(G113gat), .B(G120gat), .Z(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT31), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT31), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(KEYINPUT82), .A3(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n386_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G43gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n393_), .B(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n396_), .B(KEYINPUT83), .Z(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT1), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n415_), .A3(new_n410_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NOR4_X1   g218(.A1(KEYINPUT86), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n412_), .B2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n416_), .B(new_n419_), .C1(new_n420_), .C2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n403_), .A2(new_n404_), .B1(G155gat), .B2(G162gat), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n424_), .A2(KEYINPUT87), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT87), .B1(new_n424_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n414_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT29), .ZN(new_n429_));
  AND2_X1   g228(.A1(G197gat), .A2(G204gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT88), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G211gat), .B(G218gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT21), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n435_));
  INV_X1    g234(.A(G211gat), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n436_), .A2(G218gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(G218gat), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n437_), .A2(new_n438_), .B1(new_n431_), .B2(new_n430_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n434_), .B1(new_n440_), .B2(KEYINPUT21), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n399_), .B1(new_n429_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n399_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  AOI211_X1 g243(.A(new_n443_), .B(new_n444_), .C1(new_n428_), .C2(KEYINPUT29), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n398_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G22gat), .B(G50gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n450_), .B(KEYINPUT28), .Z(new_n451_));
  OR3_X1    g250(.A1(new_n428_), .A2(KEYINPUT29), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n428_), .B2(KEYINPUT29), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT90), .B1(new_n449_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n446_), .B(new_n447_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n414_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n424_), .A2(new_n425_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n424_), .A2(KEYINPUT87), .A3(new_n425_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n441_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n443_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n429_), .A2(new_n399_), .A3(new_n441_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n448_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT89), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n469_));
  INV_X1    g268(.A(new_n454_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n455_), .A2(new_n456_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n446_), .B(new_n448_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n474_));
  AOI211_X1 g273(.A(KEYINPUT90), .B(new_n454_), .C1(new_n467_), .C2(KEYINPUT89), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n428_), .A2(new_n389_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n389_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n480_), .B(new_n414_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(KEYINPUT4), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n428_), .A2(new_n485_), .A3(new_n389_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G29gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G85gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT0), .B(G57gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n479_), .A2(KEYINPUT4), .A3(new_n481_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n486_), .A2(new_n484_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n488_), .B(new_n493_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G190gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT26), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT26), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G190gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n365_), .A2(G183gat), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n355_), .A2(new_n501_), .A3(new_n503_), .A4(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n375_), .A2(new_n377_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n348_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n346_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .A4(new_n372_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n352_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n441_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(KEYINPUT20), .C1(new_n381_), .C2(new_n441_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G226gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT19), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT20), .B1(new_n441_), .B2(new_n510_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n381_), .A2(new_n441_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT96), .B(KEYINPUT20), .C1(new_n441_), .C2(new_n510_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n515_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G8gat), .B(G36gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G64gat), .B(G92gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT32), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n522_), .A2(KEYINPUT97), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n512_), .A2(new_n514_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n514_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT20), .B(new_n532_), .C1(new_n441_), .C2(new_n510_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n519_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n535_), .A3(new_n529_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT97), .B1(new_n522_), .B2(new_n529_), .ZN(new_n537_));
  AND4_X1   g336(.A1(new_n499_), .A2(new_n530_), .A3(new_n536_), .A4(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n498_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n533_), .B1(new_n381_), .B2(new_n441_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT21), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n542_));
  OAI221_X1 g341(.A(new_n352_), .B1(new_n542_), .B2(new_n434_), .C1(new_n368_), .C2(new_n380_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT20), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n441_), .B2(new_n510_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n532_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n527_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n531_), .A2(new_n535_), .A3(new_n528_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT92), .B(new_n527_), .C1(new_n540_), .C2(new_n546_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n539_), .A2(KEYINPUT33), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n486_), .A2(new_n483_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n496_), .B2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n482_), .A2(KEYINPUT94), .A3(new_n483_), .A4(new_n486_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n479_), .A2(new_n481_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n493_), .B1(new_n557_), .B2(new_n484_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT33), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n498_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n498_), .B2(new_n561_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n552_), .B(new_n559_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n538_), .B1(KEYINPUT95), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n550_), .A2(new_n551_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n487_), .A2(KEYINPUT33), .A3(new_n488_), .A4(new_n493_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n566_), .A2(new_n559_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n568_), .B(new_n569_), .C1(new_n563_), .C2(new_n562_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n478_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT27), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n550_), .A2(new_n572_), .A3(new_n551_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT27), .B(new_n548_), .C1(new_n522_), .C2(new_n528_), .ZN(new_n574_));
  AND4_X1   g373(.A1(new_n498_), .A2(new_n573_), .A3(new_n495_), .A4(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT98), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(new_n472_), .A3(new_n476_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n397_), .B1(new_n571_), .B2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n573_), .A2(KEYINPUT99), .A3(new_n574_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT99), .B1(new_n573_), .B2(new_n574_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n477_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(new_n396_), .A3(new_n499_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n330_), .A2(new_n331_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n590_), .A2(new_n294_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n295_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT77), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n332_), .B(new_n294_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(new_n593_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT100), .B1(new_n589_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608_));
  INV_X1    g407(.A(new_n606_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n608_), .B(new_n609_), .C1(new_n581_), .C2(new_n588_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n345_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT101), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(G1gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n499_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n202_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n612_), .A2(KEYINPUT38), .A3(new_n614_), .A4(new_n499_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n320_), .A2(new_n316_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT102), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT103), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(new_n589_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n290_), .A2(new_n609_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n344_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n499_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n616_), .A2(new_n617_), .A3(new_n628_), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n584_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G8gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n633_), .A3(G8gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n585_), .A2(G8gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n635_), .B1(new_n613_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n635_), .B(KEYINPUT40), .C1(new_n613_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1325gat));
  INV_X1    g441(.A(new_n397_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n383_), .B1(new_n625_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT41), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n612_), .A2(new_n383_), .A3(new_n643_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1326gat));
  INV_X1    g446(.A(G22gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n625_), .B2(new_n478_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT42), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n612_), .A2(new_n648_), .A3(new_n478_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n618_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n344_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n290_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT107), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n659_), .B(new_n656_), .C1(new_n607_), .C2(new_n610_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n499_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n323_), .A2(KEYINPUT43), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n589_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n577_), .A2(new_n579_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n564_), .A2(KEYINPUT95), .ZN(new_n669_));
  INV_X1    g468(.A(new_n538_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n570_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n477_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n643_), .B1(new_n668_), .B2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n667_), .B1(new_n673_), .B2(new_n587_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n581_), .A2(new_n588_), .A3(KEYINPUT105), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n323_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n319_), .A2(new_n322_), .A3(KEYINPUT106), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n675_), .A3(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n682_));
  AOI21_X1  g481(.A(new_n666_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n623_), .A2(new_n655_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n664_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n682_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n589_), .B2(new_n667_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n675_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n684_), .C1(new_n689_), .C2(new_n666_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n686_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n499_), .A2(G29gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n663_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  NOR2_X1   g492(.A1(new_n585_), .A2(G36gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n658_), .A2(new_n660_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n658_), .A2(new_n697_), .A3(new_n660_), .A4(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n686_), .A2(new_n584_), .A3(new_n690_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT46), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  AOI211_X1 g504(.A(KEYINPUT108), .B(new_n705_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1329gat));
  INV_X1    g506(.A(G43gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n396_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n691_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n661_), .B2(new_n397_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n662_), .B2(new_n478_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n478_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n691_), .B2(new_n715_), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n606_), .A2(new_n344_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n621_), .A2(new_n290_), .A3(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(G57gat), .A3(new_n499_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT110), .Z(new_n720_));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n589_), .A2(new_n609_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n290_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n724_), .A2(new_n344_), .A3(new_n324_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n627_), .B1(new_n726_), .B2(KEYINPUT109), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(KEYINPUT109), .B2(new_n726_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n720_), .B1(new_n721_), .B2(new_n728_), .ZN(G1332gat));
  INV_X1    g528(.A(G64gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n718_), .B2(new_n584_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n726_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n730_), .A3(new_n584_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n718_), .B2(new_n643_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n737_), .A3(new_n643_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n718_), .A2(new_n478_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G78gat), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n477_), .A2(G78gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n726_), .B2(new_n746_), .ZN(G1335gat));
  NAND3_X1  g546(.A1(new_n290_), .A2(new_n344_), .A3(new_n619_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n722_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n499_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n681_), .A2(new_n682_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n666_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n724_), .A2(new_n606_), .A3(new_n655_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n627_), .A2(new_n239_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n750_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n749_), .A2(new_n240_), .A3(new_n584_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n755_), .A2(new_n584_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n240_), .ZN(G1337gat));
  NAND2_X1  g559(.A1(new_n755_), .A2(new_n643_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n204_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n396_), .A2(new_n762_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n761_), .A2(G99gat), .B1(new_n749_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n749_), .A2(new_n205_), .A3(new_n478_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n753_), .A2(new_n478_), .A3(new_n754_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(G106gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g572(.A1(new_n287_), .A2(new_n289_), .A3(new_n717_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n287_), .A2(new_n289_), .A3(KEYINPUT114), .A4(new_n717_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n323_), .A3(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n776_), .A2(new_n323_), .A3(new_n777_), .A4(new_n779_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n606_), .A2(new_n284_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n272_), .A2(new_n786_), .A3(new_n263_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n262_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n273_), .A2(new_n786_), .A3(new_n277_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n282_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT56), .B(new_n282_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n785_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n591_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n603_), .C1(new_n597_), .C2(new_n595_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n605_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n288_), .B2(new_n284_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT57), .B(new_n654_), .C1(new_n798_), .C2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n284_), .A2(new_n605_), .A3(new_n800_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n324_), .B1(new_n805_), .B2(KEYINPUT58), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n807_), .B(new_n804_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n803_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n785_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n789_), .A2(new_n790_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n282_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n797_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n810_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n802_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n619_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n344_), .B1(new_n809_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n784_), .A2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n586_), .A2(new_n396_), .A3(new_n627_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT117), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n654_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n815_), .A2(new_n816_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n807_), .B1(new_n832_), .B2(new_n804_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n805_), .A2(KEYINPUT58), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n324_), .A3(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n827_), .A2(new_n831_), .A3(new_n803_), .A4(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n344_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n784_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(new_n823_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n826_), .B1(new_n839_), .B2(new_n824_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n609_), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n842_), .A3(new_n606_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1340gat));
  OAI21_X1  g643(.A(G120gat), .B1(new_n840_), .B2(new_n724_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  AOI21_X1  g645(.A(G120gat), .B1(new_n290_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT118), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n846_), .B2(G120gat), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n839_), .B(new_n848_), .C1(new_n847_), .C2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n845_), .A2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n839_), .B2(new_n655_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n840_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n655_), .A2(G127gat), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT119), .Z(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n854_), .B2(new_n856_), .ZN(G1342gat));
  OAI21_X1  g656(.A(G134gat), .B1(new_n840_), .B2(new_n323_), .ZN(new_n858_));
  INV_X1    g657(.A(G134gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n620_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n839_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(G1343gat));
  AOI21_X1  g661(.A(new_n783_), .B1(new_n836_), .B2(new_n344_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n397_), .A2(new_n478_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(new_n627_), .A3(new_n584_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT120), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n829_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n809_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n655_), .B1(new_n870_), .B2(new_n831_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n868_), .B(new_n865_), .C1(new_n871_), .C2(new_n783_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n606_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n290_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n655_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n873_), .B2(new_n680_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n860_), .A2(new_n881_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n867_), .B2(new_n872_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT121), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n873_), .A2(new_n881_), .A3(new_n860_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n679_), .B1(new_n867_), .B2(new_n872_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n886_), .B(new_n887_), .C1(new_n881_), .C2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n889_), .ZN(G1347gat));
  XNOR2_X1  g689(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n585_), .A2(new_n499_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n822_), .A2(new_n643_), .A3(new_n477_), .A4(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n609_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT22), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G169gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n370_), .B1(new_n894_), .B2(new_n891_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n896_), .B2(new_n898_), .ZN(G1348gat));
  NAND2_X1  g698(.A1(new_n838_), .A2(new_n477_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n892_), .A2(new_n643_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n900_), .A2(new_n371_), .A3(new_n724_), .A4(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n371_), .B1(new_n893_), .B2(new_n724_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n903_), .A2(KEYINPUT123), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(KEYINPUT123), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  AOI211_X1 g705(.A(new_n344_), .B(new_n893_), .C1(new_n355_), .C2(new_n504_), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n900_), .A2(new_n344_), .A3(new_n901_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n354_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n893_), .B2(new_n323_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n860_), .A2(new_n353_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n893_), .B2(new_n911_), .ZN(G1351gat));
  XOR2_X1   g711(.A(KEYINPUT124), .B(G197gat), .Z(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n864_), .A2(new_n499_), .A3(new_n585_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n838_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n609_), .ZN(new_n917_));
  MUX2_X1   g716(.A(new_n913_), .B(new_n914_), .S(new_n917_), .Z(G1352gat));
  INV_X1    g717(.A(new_n916_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n290_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g720(.A1(new_n916_), .A2(new_n344_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT63), .B(G211gat), .Z(new_n923_));
  AOI21_X1  g722(.A(KEYINPUT125), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n923_), .ZN(new_n925_));
  OR2_X1    g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n922_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n927_), .B2(KEYINPUT125), .ZN(G1354gat));
  NAND2_X1  g727(.A1(new_n324_), .A2(G218gat), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT126), .Z(new_n930_));
  NAND2_X1  g729(.A1(new_n919_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n916_), .A2(new_n620_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(G218gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT127), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n931_), .B(new_n935_), .C1(new_n932_), .C2(G218gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(G1355gat));
endmodule


