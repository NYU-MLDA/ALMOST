//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n203_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT78), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT77), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT77), .B1(new_n215_), .B2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OAI221_X1 g016(.A(new_n208_), .B1(new_n209_), .B2(new_n211_), .C1(new_n213_), .C2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n220_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT79), .B(G176gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n211_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n218_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT30), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(G15gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G43gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G99gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  NAND3_X1  g034(.A1(new_n228_), .A2(new_n229_), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n229_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n236_), .B(KEYINPUT83), .C1(new_n228_), .C2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n239_), .A2(new_n240_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT82), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT31), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n238_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n238_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT3), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(KEYINPUT2), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n258_), .A2(new_n259_), .B1(new_n256_), .B2(KEYINPUT2), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n255_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT86), .Z(new_n263_));
  OAI211_X1 g062(.A(new_n252_), .B(new_n253_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n252_), .A2(KEYINPUT1), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(G155gat), .A3(G162gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n265_), .A2(new_n267_), .A3(new_n253_), .A4(KEYINPUT84), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n258_), .A2(new_n259_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(new_n254_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n268_), .B(new_n270_), .C1(KEYINPUT84), .C2(new_n267_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n264_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n272_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G22gat), .B(G50gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G78gat), .B(G106gat), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  INV_X1    g082(.A(G204gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT90), .B1(new_n284_), .B2(G197gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(KEYINPUT21), .A3(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G197gat), .B(G204gat), .Z(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n286_), .B(new_n287_), .C1(KEYINPUT21), .C2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT89), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n293_));
  INV_X1    g092(.A(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(G228gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(G228gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n293_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT91), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n280_), .A2(new_n282_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n282_), .B1(new_n280_), .B2(new_n300_), .ZN(new_n302_));
  OAI22_X1  g101(.A1(new_n301_), .A2(new_n302_), .B1(KEYINPUT91), .B2(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n280_), .A2(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n281_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n299_), .A2(KEYINPUT91), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n280_), .A2(new_n282_), .A3(new_n300_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n227_), .A2(new_n290_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n225_), .A2(new_n219_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT92), .ZN(new_n313_));
  INV_X1    g112(.A(new_n209_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n212_), .A2(new_n214_), .B1(new_n314_), .B2(new_n210_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n208_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(KEYINPUT20), .B(new_n311_), .C1(new_n317_), .C2(new_n291_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT19), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n227_), .A2(new_n290_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n291_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT94), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n318_), .A2(new_n320_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n333_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n244_), .A2(new_n241_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n272_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n246_), .B2(new_n272_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT95), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n272_), .A2(new_n246_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(KEYINPUT4), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n340_), .B2(KEYINPUT4), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n344_), .B(new_n348_), .C1(new_n351_), .C2(new_n343_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n334_), .A2(new_n337_), .A3(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n341_), .A2(new_n343_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n343_), .B2(new_n351_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(new_n348_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT33), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n355_), .A2(KEYINPUT33), .A3(new_n348_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n312_), .A2(new_n316_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT20), .B1(new_n361_), .B2(new_n290_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n320_), .B1(new_n322_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n336_), .A2(KEYINPUT32), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n365_), .B2(new_n327_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n355_), .A2(new_n348_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n357_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n310_), .B1(new_n360_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n357_), .A2(new_n368_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n334_), .A2(new_n337_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n364_), .A2(new_n333_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n373_), .A2(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n309_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n251_), .B1(new_n370_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n308_), .A3(new_n303_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n377_), .A2(new_n303_), .A3(KEYINPUT96), .A4(new_n308_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n382_), .A2(new_n372_), .A3(new_n251_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT97), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n250_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n387_), .A2(KEYINPUT97), .A3(new_n372_), .A4(new_n383_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n379_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G15gat), .B(G22gat), .ZN(new_n390_));
  INV_X1    g189(.A(G1gat), .ZN(new_n391_));
  INV_X1    g190(.A(G8gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT14), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G8gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  XNOR2_X1  g195(.A(G57gat), .B(G64gat), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT11), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(KEYINPUT11), .ZN(new_n399_));
  XOR2_X1   g198(.A(G71gat), .B(G78gat), .Z(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n399_), .A2(new_n400_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n396_), .B(new_n403_), .Z(new_n404_));
  NAND2_X1  g203(.A1(G231gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G127gat), .B(G155gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G183gat), .B(G211gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT17), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n411_), .A2(KEYINPUT17), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G190gat), .B(G218gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT71), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G134gat), .B(G162gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT36), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT10), .B(G99gat), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT64), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(KEYINPUT64), .ZN(new_n424_));
  AOI21_X1  g223(.A(G106gat), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G85gat), .B(G92gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT9), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G99gat), .A2(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT6), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT9), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(G85gat), .A3(G92gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n427_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n425_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438_));
  INV_X1    g237(.A(G99gat), .ZN(new_n439_));
  INV_X1    g238(.A(G106gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT7), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT7), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n443_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n432_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT8), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n426_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n445_), .B2(new_n426_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n426_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT67), .B1(new_n453_), .B2(new_n447_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n437_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n450_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(KEYINPUT67), .A3(new_n447_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT68), .A3(new_n437_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n457_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n436_), .B1(new_n453_), .B2(new_n447_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G232gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT34), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n469_), .A2(new_n465_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n468_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n470_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n475_), .A2(new_n476_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n421_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n420_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n483_), .A3(new_n477_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT72), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n389_), .A2(new_n416_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n469_), .A2(new_n403_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n469_), .A2(new_n403_), .ZN(new_n494_));
  OR3_X1    g293(.A1(new_n493_), .A2(KEYINPUT66), .A3(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n493_), .B2(KEYINPUT66), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n401_), .A2(KEYINPUT12), .A3(new_n402_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT68), .B1(new_n460_), .B2(new_n437_), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n456_), .B(new_n436_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n494_), .A2(KEYINPUT12), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n496_), .B1(new_n469_), .B2(new_n403_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n498_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G120gat), .B(G148gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT5), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G176gat), .B(G204gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n511_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n498_), .A2(new_n506_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n512_), .A2(KEYINPUT13), .A3(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT69), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n465_), .B(KEYINPUT75), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n396_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT76), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n523_), .A2(new_n396_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n396_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n467_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n522_), .B2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G113gat), .B(G141gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(G169gat), .B(G197gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n531_), .B(new_n534_), .Z(new_n535_));
  NOR2_X1   g334(.A1(new_n521_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n491_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n537_), .B(KEYINPUT98), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n391_), .A3(new_n371_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT38), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n389_), .A2(new_n535_), .A3(new_n519_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n486_), .A2(new_n416_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n391_), .B1(new_n544_), .B2(new_n371_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n540_), .B2(new_n539_), .ZN(G1324gat));
  INV_X1    g346(.A(KEYINPUT39), .ZN(new_n548_));
  OAI21_X1  g347(.A(G8gat), .B1(new_n548_), .B2(KEYINPUT99), .ZN(new_n549_));
  INV_X1    g348(.A(new_n377_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(KEYINPUT99), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n377_), .A2(G8gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(new_n538_), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT40), .ZN(G1325gat));
  AOI21_X1  g355(.A(new_n231_), .B1(new_n544_), .B2(new_n251_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT41), .ZN(new_n558_));
  INV_X1    g357(.A(new_n537_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n231_), .A3(new_n251_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(G1326gat));
  INV_X1    g360(.A(G22gat), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n544_), .B2(new_n309_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT42), .Z(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n562_), .A3(new_n309_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(G1327gat));
  INV_X1    g365(.A(new_n416_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n485_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n542_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G29gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n371_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT101), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n386_), .A2(new_n388_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n379_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT43), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n490_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT43), .B1(new_n389_), .B2(new_n489_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT100), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n519_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n535_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n416_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT100), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT44), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT44), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n586_), .A3(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n371_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n572_), .B1(new_n589_), .B2(G29gat), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT101), .B(new_n570_), .C1(new_n588_), .C2(new_n371_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n571_), .B1(new_n590_), .B2(new_n591_), .ZN(G1328gat));
  INV_X1    g391(.A(KEYINPUT104), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT46), .ZN(new_n594_));
  INV_X1    g393(.A(G36gat), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n542_), .A2(new_n595_), .A3(new_n550_), .A4(new_n568_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n579_), .A2(new_n586_), .A3(new_n583_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n586_), .B1(new_n579_), .B2(new_n583_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n550_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n601_), .B2(G36gat), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT103), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n594_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT103), .B(new_n598_), .C1(new_n601_), .C2(G36gat), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n593_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n598_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n377_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(new_n595_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT103), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n602_), .A2(new_n603_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT104), .A4(new_n594_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n602_), .A2(KEYINPUT46), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n606_), .A2(new_n612_), .A3(new_n613_), .ZN(G1329gat));
  AOI21_X1  g413(.A(G43gat), .B1(new_n569_), .B2(new_n251_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n251_), .A2(G43gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n588_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g418(.A(G50gat), .B1(new_n569_), .B2(new_n309_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n309_), .A2(G50gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n588_), .B2(new_n621_), .ZN(G1331gat));
  NOR2_X1   g421(.A1(new_n580_), .A2(new_n581_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n491_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(G57gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n371_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n389_), .A2(new_n581_), .A3(new_n520_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n543_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G57gat), .B1(new_n628_), .B2(new_n372_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(G1332gat));
  OAI21_X1  g429(.A(G64gat), .B1(new_n628_), .B2(new_n377_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(G64gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n624_), .A2(new_n634_), .A3(new_n550_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1333gat));
  OAI21_X1  g435(.A(G71gat), .B1(new_n628_), .B2(new_n250_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(G71gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n624_), .A2(new_n640_), .A3(new_n251_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1334gat));
  OAI21_X1  g441(.A(G78gat), .B1(new_n628_), .B2(new_n310_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT50), .ZN(new_n644_));
  INV_X1    g443(.A(G78gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n624_), .A2(new_n645_), .A3(new_n309_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1335gat));
  NAND2_X1  g446(.A1(new_n577_), .A2(new_n578_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n580_), .A2(new_n567_), .A3(new_n581_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(G85gat), .A3(new_n371_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n627_), .A2(new_n568_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G85gat), .B1(new_n653_), .B2(new_n371_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(KEYINPUT107), .B2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(KEYINPUT107), .B2(new_n654_), .ZN(G1336gat));
  NAND3_X1  g455(.A1(new_n651_), .A2(G92gat), .A3(new_n550_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  AOI21_X1  g457(.A(G92gat), .B1(new_n653_), .B2(new_n550_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n658_), .B2(new_n659_), .ZN(G1337gat));
  INV_X1    g460(.A(KEYINPUT111), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n423_), .A2(new_n424_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n653_), .A2(new_n251_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n651_), .A2(new_n251_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n650_), .A2(new_n250_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n439_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n665_), .B1(new_n667_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT51), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n662_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT109), .B1(new_n666_), .B2(G99gat), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n669_), .A2(new_n668_), .A3(new_n439_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n664_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT110), .B1(new_n676_), .B2(KEYINPUT51), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT110), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n671_), .A2(new_n679_), .A3(new_n672_), .ZN(new_n680_));
  OAI22_X1  g479(.A1(new_n673_), .A2(new_n677_), .B1(new_n678_), .B2(new_n680_), .ZN(G1338gat));
  NAND3_X1  g480(.A1(new_n653_), .A2(new_n440_), .A3(new_n309_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT52), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n651_), .A2(new_n309_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(G106gat), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT52), .B(new_n440_), .C1(new_n651_), .C2(new_n309_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g487(.A1(new_n387_), .A2(new_n383_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n371_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n503_), .A2(new_n504_), .A3(new_n492_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n506_), .A2(KEYINPUT55), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT55), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n503_), .A2(new_n504_), .A3(new_n693_), .A4(new_n505_), .ZN(new_n694_));
  AOI221_X4 g493(.A(KEYINPUT113), .B1(new_n691_), .B2(new_n496_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n692_), .A2(new_n694_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n691_), .A2(new_n496_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n511_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT114), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT56), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n703_), .A2(new_n581_), .A3(new_n514_), .A4(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n530_), .A2(G229gat), .A3(G233gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n525_), .A2(new_n526_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n534_), .B1(new_n707_), .B2(new_n522_), .ZN(new_n708_));
  AOI22_X1  g507(.A1(new_n531_), .A2(new_n534_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n515_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT115), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n486_), .B1(new_n705_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT57), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT56), .B(new_n511_), .C1(new_n695_), .C2(new_n699_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT116), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n494_), .A2(KEYINPUT12), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n462_), .B2(new_n500_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n693_), .B1(new_n718_), .B2(new_n505_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n694_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n698_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT113), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n697_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT56), .B1(new_n724_), .B2(new_n511_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n716_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT116), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n700_), .A2(new_n727_), .A3(new_n702_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n709_), .A2(new_n514_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT117), .B1(new_n726_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT58), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n700_), .A2(new_n702_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(KEYINPUT116), .A3(new_n715_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT117), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n732_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(KEYINPUT118), .A3(new_n490_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n734_), .A2(KEYINPUT58), .A3(new_n728_), .A4(new_n729_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT118), .B1(new_n737_), .B2(new_n490_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n714_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT119), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT119), .B(new_n714_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n416_), .A3(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n489_), .A2(new_n567_), .A3(new_n535_), .A4(new_n580_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n690_), .B1(new_n746_), .B2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G113gat), .B1(new_n751_), .B2(new_n581_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n746_), .A2(new_n750_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n690_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT59), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT59), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n742_), .A2(new_n416_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n757_), .B(new_n754_), .C1(new_n758_), .C2(new_n749_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n756_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n581_), .B2(KEYINPUT120), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(KEYINPUT120), .B2(new_n761_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n752_), .B1(new_n760_), .B2(new_n763_), .ZN(G1340gat));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n521_), .A3(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G120gat), .ZN(new_n766_));
  INV_X1    g565(.A(G120gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n580_), .B2(KEYINPUT60), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n751_), .B(new_n768_), .C1(KEYINPUT60), .C2(new_n767_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1341gat));
  NAND3_X1  g569(.A1(new_n756_), .A2(new_n567_), .A3(new_n759_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G127gat), .ZN(new_n772_));
  OR3_X1    g571(.A1(new_n755_), .A2(G127gat), .A3(new_n416_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1342gat));
  NAND3_X1  g573(.A1(new_n753_), .A2(new_n486_), .A3(new_n754_), .ZN(new_n775_));
  INV_X1    g574(.A(G134gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n489_), .A2(new_n776_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n759_), .B(new_n778_), .C1(new_n751_), .C2(new_n757_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n777_), .A2(new_n779_), .A3(KEYINPUT121), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1343gat));
  NOR3_X1   g583(.A1(new_n310_), .A2(new_n372_), .A3(new_n251_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n753_), .A2(new_n377_), .A3(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n535_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT122), .B(G141gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1344gat));
  NOR2_X1   g588(.A1(new_n786_), .A2(new_n520_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT123), .B(G148gat), .Z(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1345gat));
  NOR2_X1   g591(.A1(new_n786_), .A2(new_n416_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT61), .B(G155gat), .Z(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1346gat));
  OAI21_X1  g594(.A(G162gat), .B1(new_n786_), .B2(new_n489_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n485_), .A2(G162gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n786_), .B2(new_n797_), .ZN(G1347gat));
  NOR2_X1   g597(.A1(new_n758_), .A2(new_n749_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n550_), .A2(new_n372_), .A3(new_n251_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n310_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n799_), .A2(new_n535_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT62), .ZN(new_n804_));
  OR3_X1    g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n205_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(new_n205_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n224_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(G1348gat));
  NOR3_X1   g607(.A1(new_n799_), .A2(new_n580_), .A3(new_n802_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n223_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n800_), .A2(new_n206_), .ZN(new_n812_));
  AND4_X1   g611(.A1(new_n310_), .A2(new_n753_), .A3(new_n521_), .A4(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT124), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n567_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n749_), .B1(new_n815_), .B2(new_n745_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n309_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n521_), .A3(new_n812_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n818_), .B(new_n819_), .C1(new_n810_), .C2(new_n809_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n814_), .A2(new_n820_), .ZN(G1349gat));
  NAND3_X1  g620(.A1(new_n817_), .A2(new_n567_), .A3(new_n801_), .ZN(new_n822_));
  INV_X1    g621(.A(G183gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n799_), .A2(new_n802_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n416_), .A2(new_n214_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n822_), .A2(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(G1350gat));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n212_), .A3(new_n486_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n490_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n828_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT125), .B1(new_n828_), .B2(G190gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(G1351gat));
  NAND2_X1  g630(.A1(new_n309_), .A2(new_n372_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(new_n377_), .A3(new_n251_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n753_), .A2(KEYINPUT126), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT126), .ZN(new_n835_));
  INV_X1    g634(.A(new_n833_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n816_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G197gat), .B1(new_n838_), .B2(new_n581_), .ZN(new_n839_));
  INV_X1    g638(.A(G197gat), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n840_), .B(new_n535_), .C1(new_n834_), .C2(new_n837_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1352gat));
  NOR2_X1   g641(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n520_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n838_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n845_), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n847_), .B(new_n843_), .C1(new_n834_), .C2(new_n837_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1353gat));
  OR2_X1    g648(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n838_), .B2(new_n567_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT63), .B(G211gat), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n416_), .B(new_n852_), .C1(new_n834_), .C2(new_n837_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1354gat));
  INV_X1    g653(.A(G218gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n838_), .A2(new_n855_), .A3(new_n486_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n489_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n855_), .B2(new_n857_), .ZN(G1355gat));
endmodule


