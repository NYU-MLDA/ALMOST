//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT91), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT90), .B(G197gat), .ZN(new_n206_));
  AOI22_X1  g005(.A1(new_n205_), .A2(G197gat), .B1(new_n206_), .B2(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT91), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G204gat), .ZN(new_n214_));
  INV_X1    g013(.A(G197gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n217_), .A2(new_n218_), .A3(G204gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT21), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(G204gat), .B1(new_n217_), .B2(new_n218_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(new_n208_), .C1(new_n215_), .C2(new_n204_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n209_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT92), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n220_), .A2(KEYINPUT92), .A3(new_n209_), .A4(new_n222_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n210_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT26), .B(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT82), .ZN(new_n231_));
  AND2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT23), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(G183gat), .A3(G190gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n234_), .A2(KEYINPUT24), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n233_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n228_), .A2(new_n229_), .A3(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n231_), .A2(new_n239_), .A3(new_n241_), .A4(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n238_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n232_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT22), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT22), .B1(new_n249_), .B2(new_n250_), .ZN(new_n252_));
  INV_X1    g051(.A(G176gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n248_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n244_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT20), .B1(new_n227_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n234_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n233_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n245_), .A4(new_n230_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT22), .B(G169gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n253_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n248_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  AOI211_X1 g066(.A(new_n210_), .B(new_n267_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n203_), .B1(new_n258_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n225_), .A2(new_n226_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n210_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n267_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n203_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n227_), .A2(new_n257_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n273_), .A2(KEYINPUT20), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT32), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n267_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT20), .B1(new_n227_), .B2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n270_), .A2(new_n257_), .A3(new_n271_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n203_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n272_), .A2(new_n256_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n227_), .A2(new_n286_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(KEYINPUT20), .A3(new_n274_), .A4(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n289_), .A2(new_n292_), .A3(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT87), .B1(new_n297_), .B2(KEYINPUT1), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(G155gat), .A4(G162gat), .ZN(new_n301_));
  INV_X1    g100(.A(G155gat), .ZN(new_n302_));
  INV_X1    g101(.A(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(KEYINPUT1), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n298_), .A2(new_n301_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(G141gat), .ZN(new_n308_));
  INV_X1    g107(.A(G148gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .A4(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT88), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n304_), .A2(new_n297_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n311_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT97), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n318_), .A2(new_n320_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT88), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n311_), .A3(new_n327_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n296_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n333_), .B2(new_n311_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT4), .B1(new_n336_), .B2(new_n324_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n295_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n334_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(new_n336_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n294_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343_));
  INV_X1    g142(.A(G85gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n285_), .B(new_n293_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n352_), .A2(KEYINPUT33), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n338_), .A2(new_n341_), .A3(new_n347_), .A4(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n352_), .B1(KEYINPUT99), .B2(KEYINPUT33), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n282_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n272_), .B2(new_n267_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n274_), .B1(new_n359_), .B2(new_n275_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n258_), .A2(new_n268_), .A3(new_n203_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n289_), .A2(new_n292_), .A3(new_n282_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n294_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n340_), .A2(new_n295_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n348_), .A3(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n356_), .A2(new_n362_), .A3(new_n363_), .A4(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n342_), .A2(new_n348_), .A3(new_n355_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n351_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(G50gat), .B1(new_n323_), .B2(KEYINPUT29), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT28), .B(G22gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  INV_X1    g171(.A(G50gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n333_), .A2(new_n372_), .A3(new_n373_), .A4(new_n311_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n371_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT94), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n375_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n323_), .A2(KEYINPUT29), .ZN(new_n382_));
  AND2_X1   g181(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(G228gat), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT93), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n272_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n272_), .A2(new_n382_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n385_), .B(KEYINPUT93), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n378_), .A2(new_n381_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n379_), .A2(new_n375_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n388_), .A2(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n387_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(KEYINPUT94), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n369_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n369_), .A2(new_n401_), .A3(KEYINPUT100), .ZN(new_n405_));
  INV_X1    g204(.A(new_n400_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n397_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n349_), .A2(new_n350_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n289_), .A2(new_n292_), .A3(new_n282_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n282_), .B1(new_n269_), .B2(new_n276_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT101), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT101), .B1(new_n277_), .B2(new_n357_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n362_), .A2(new_n410_), .A3(new_n363_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n408_), .B(new_n409_), .C1(new_n416_), .C2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n404_), .A2(new_n405_), .A3(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n256_), .B(KEYINPUT30), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G71gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(new_n328_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT85), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G43gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G99gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n427_), .B(new_n429_), .Z(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n422_), .B(new_n327_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT86), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT102), .B1(new_n416_), .B2(new_n418_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT102), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n277_), .A2(new_n357_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n363_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n440_), .B2(KEYINPUT101), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n438_), .B(new_n417_), .C1(new_n441_), .C2(new_n410_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n408_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n409_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n435_), .A2(new_n444_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n420_), .A2(new_n436_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G29gat), .B(G36gat), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(G50gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT72), .B(G43gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(G50gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT15), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n447_), .B(G50gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n449_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT15), .B1(new_n458_), .B2(new_n451_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n461_));
  INV_X1    g260(.A(G99gat), .ZN(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n467_));
  OAI22_X1  g266(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G85gat), .A2(G92gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n469_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT8), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT68), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT9), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT64), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n471_), .A2(new_n481_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT64), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n473_), .A2(new_n483_), .A3(new_n478_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n480_), .A2(new_n482_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT10), .B(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n463_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n486_), .A2(new_n489_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n477_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n475_), .A2(KEYINPUT68), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n469_), .A2(new_n493_), .A3(new_n474_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(KEYINPUT8), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n460_), .A2(new_n496_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n458_), .A2(new_n451_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(new_n505_), .A3(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n502_), .A2(new_n497_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n503_), .A2(new_n510_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G190gat), .B(G218gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(new_n303_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT73), .B(G134gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n509_), .A2(KEYINPUT36), .A3(new_n511_), .A4(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(KEYINPUT36), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n509_), .A2(new_n511_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI211_X1 g321(.A(KEYINPUT74), .B(new_n518_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT104), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n446_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT105), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT13), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G71gat), .B(G78gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(G57gat), .A2(G64gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT11), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G57gat), .A2(G64gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT11), .B1(new_n537_), .B2(new_n532_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n531_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n530_), .B(KEYINPUT11), .C1(new_n532_), .C2(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n495_), .A2(new_n477_), .A3(new_n490_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n541_), .B(KEYINPUT69), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n492_), .A2(KEYINPUT8), .A3(new_n494_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n477_), .A2(new_n490_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n548_), .B(KEYINPUT12), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n541_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT12), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT71), .B1(new_n547_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n542_), .A2(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT70), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n552_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n544_), .B1(new_n563_), .B2(new_n542_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G204gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT5), .B(G176gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n562_), .A2(new_n565_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n529_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(KEYINPUT13), .A3(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n505_), .A2(new_n453_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G8gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT76), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582_));
  INV_X1    g381(.A(G1gat), .ZN(new_n583_));
  INV_X1    g382(.A(G8gat), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT14), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n580_), .A2(KEYINPUT76), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n580_), .A2(KEYINPUT76), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n585_), .A3(new_n582_), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n458_), .A2(KEYINPUT15), .A3(new_n451_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n579_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n505_), .A2(new_n591_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n505_), .A2(new_n591_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n505_), .A2(new_n591_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n308_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT79), .B(G113gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n597_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT80), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT81), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n608_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n610_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT81), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(new_n602_), .A3(new_n607_), .A4(new_n612_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n578_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n591_), .B(KEYINPUT77), .Z(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(new_n548_), .Z(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n624_), .A2(new_n541_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n541_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .A4(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n621_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT103), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n528_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n409_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n524_), .A2(KEYINPUT37), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n524_), .A2(KEYINPUT37), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n640_), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n446_), .A2(new_n620_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n583_), .A3(new_n444_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT38), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n650_), .ZN(G1324gat));
  AND2_X1   g450(.A1(new_n437_), .A2(new_n442_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n584_), .A3(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n528_), .A2(new_n652_), .A3(new_n642_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(G8gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n654_), .B2(G8gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1325gat));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n436_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G15gat), .B1(new_n643_), .B2(new_n436_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n667_), .B(G15gat), .C1(new_n643_), .C2(new_n436_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n663_), .B1(new_n669_), .B2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n648_), .A2(new_n672_), .A3(new_n408_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n528_), .A2(new_n408_), .A3(new_n642_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G22gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1327gat));
  NOR2_X1   g479(.A1(new_n620_), .A2(new_n640_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n420_), .A2(new_n436_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n443_), .A2(new_n445_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n645_), .A2(new_n646_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n686_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n446_), .A2(KEYINPUT43), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n681_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n681_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n409_), .ZN(new_n695_));
  INV_X1    g494(.A(G29gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n681_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n526_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n446_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n444_), .A2(new_n696_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT108), .B1(new_n697_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  OAI221_X1 g504(.A(new_n705_), .B1(new_n701_), .B2(new_n702_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1328gat));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n708_), .A3(new_n652_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT45), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n700_), .A2(new_n711_), .A3(new_n708_), .A4(new_n652_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(KEYINPUT110), .A3(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n692_), .A2(KEYINPUT109), .A3(new_n652_), .A4(new_n693_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n692_), .A2(new_n652_), .A3(new_n693_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT46), .B(new_n713_), .C1(new_n715_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n718_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n722_), .A2(KEYINPUT110), .A3(G36gat), .A4(new_n714_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n713_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n720_), .A2(new_n725_), .ZN(G1329gat));
  INV_X1    g525(.A(new_n435_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G43gat), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n701_), .A2(new_n436_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n694_), .A2(new_n728_), .B1(G43gat), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n694_), .B2(new_n401_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n700_), .A2(new_n373_), .A3(new_n408_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1331gat));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n446_), .A2(new_n647_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n578_), .A2(new_n619_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n738_), .B2(new_n409_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT111), .Z(new_n740_));
  AND3_X1   g539(.A1(new_n528_), .A2(new_n640_), .A3(new_n737_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n409_), .A2(new_n735_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(G1332gat));
  INV_X1    g542(.A(new_n738_), .ZN(new_n744_));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n652_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n652_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G64gat), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1333gat));
  OR3_X1    g550(.A1(new_n738_), .A2(G71gat), .A3(new_n436_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n741_), .A2(new_n662_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G71gat), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT49), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT49), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1334gat));
  OR3_X1    g556(.A1(new_n738_), .A2(G78gat), .A3(new_n401_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n528_), .A2(new_n408_), .A3(new_n640_), .A4(new_n737_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G78gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G78gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT112), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n758_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1335gat));
  NOR3_X1   g566(.A1(new_n578_), .A2(new_n619_), .A3(new_n640_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n685_), .A2(new_n526_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n444_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n687_), .A2(new_n689_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n768_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n409_), .A2(new_n344_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1336gat));
  AOI21_X1  g574(.A(G92gat), .B1(new_n769_), .B2(new_n652_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n652_), .A2(G92gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(G1337gat));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779_));
  OAI21_X1  g578(.A(G99gat), .B1(new_n772_), .B2(new_n436_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n769_), .A2(new_n488_), .A3(new_n727_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n782_), .A2(new_n785_), .A3(new_n783_), .A4(new_n779_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1338gat));
  OAI21_X1  g588(.A(G106gat), .B1(new_n772_), .B2(new_n401_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT52), .B(G106gat), .C1(new_n772_), .C2(new_n401_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n769_), .A2(new_n463_), .A3(new_n408_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT115), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n796_), .B(new_n798_), .ZN(G1339gat));
  NAND3_X1  g598(.A1(new_n594_), .A2(new_n598_), .A3(new_n596_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n595_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n607_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n609_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n554_), .B2(new_n561_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n555_), .A2(new_n559_), .A3(KEYINPUT55), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n551_), .B(new_n542_), .C1(new_n552_), .C2(KEYINPUT12), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  INV_X1    g606(.A(new_n544_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n569_), .B1(new_n804_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT56), .B(new_n569_), .C1(new_n804_), .C2(new_n811_), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n572_), .B(new_n803_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT58), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n803_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n571_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT121), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n822_), .A3(new_n686_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n803_), .B1(new_n575_), .B2(new_n571_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n812_), .A2(KEYINPUT119), .A3(new_n813_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n826_), .A2(new_n571_), .A3(new_n619_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n814_), .A2(new_n828_), .A3(new_n815_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n825_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n824_), .B1(new_n830_), .B2(new_n526_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n619_), .A2(new_n571_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n826_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n825_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n526_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n823_), .A2(new_n831_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n639_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n647_), .A2(new_n577_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  INV_X1    g639(.A(new_n619_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT54), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n839_), .A2(KEYINPUT117), .A3(new_n840_), .A4(new_n841_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n838_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n443_), .A2(new_n444_), .A3(new_n727_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n835_), .B2(KEYINPUT57), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT120), .B(new_n824_), .C1(new_n830_), .C2(new_n526_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n823_), .A4(new_n836_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n639_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n850_), .B1(new_n857_), .B2(new_n848_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n619_), .B(new_n852_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G113gat), .ZN(new_n861_));
  INV_X1    g660(.A(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(new_n862_), .A3(new_n619_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(KEYINPUT122), .A3(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1340gat));
  NAND2_X1  g667(.A1(new_n857_), .A2(new_n848_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n850_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT60), .B1(new_n577_), .B2(new_n872_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n871_), .A2(KEYINPUT60), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n852_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n873_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n876_), .A2(new_n578_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n874_), .B1(new_n878_), .B2(new_n872_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n858_), .B2(new_n640_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n876_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n640_), .A2(G127gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1342gat));
  AOI21_X1  g682(.A(G134gat), .B1(new_n858_), .B2(new_n526_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n686_), .A2(G134gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n881_), .B2(new_n885_), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n662_), .A2(new_n401_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n888_), .A2(new_n409_), .A3(new_n652_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n869_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n841_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n308_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n578_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n309_), .ZN(G1345gat));
  AND2_X1   g693(.A1(new_n869_), .A2(new_n889_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n302_), .A3(new_n640_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G155gat), .B1(new_n890_), .B2(new_n639_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n899_), .A3(new_n897_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  AOI21_X1  g702(.A(new_n303_), .B1(new_n895_), .B2(new_n686_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n890_), .A2(G162gat), .A3(new_n699_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n904_), .A2(new_n905_), .A3(KEYINPUT124), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n895_), .A2(new_n303_), .A3(new_n526_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G162gat), .B1(new_n890_), .B2(new_n688_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n906_), .A2(new_n910_), .ZN(G1347gat));
  INV_X1    g710(.A(new_n849_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n652_), .A2(new_n409_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n662_), .ZN(new_n914_));
  OR3_X1    g713(.A1(new_n914_), .A2(KEYINPUT125), .A3(new_n841_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT125), .B1(new_n914_), .B2(new_n841_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n401_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n912_), .B2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT62), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n914_), .A2(new_n408_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n849_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n264_), .A3(new_n619_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n923_), .ZN(G1348gat));
  NAND3_X1  g723(.A1(new_n922_), .A2(new_n253_), .A3(new_n577_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n869_), .A2(new_n577_), .A3(new_n920_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n253_), .B2(new_n926_), .ZN(G1349gat));
  NOR2_X1   g726(.A1(new_n921_), .A2(new_n639_), .ZN(new_n928_));
  MUX2_X1   g727(.A(G183gat), .B(new_n228_), .S(new_n928_), .Z(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n921_), .B2(new_n688_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n526_), .A2(new_n229_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n921_), .B2(new_n931_), .ZN(G1351gat));
  AOI21_X1  g731(.A(new_n888_), .B1(new_n857_), .B2(new_n848_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n913_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n841_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n215_), .ZN(G1352gat));
  OAI21_X1  g735(.A(G204gat), .B1(new_n934_), .B2(new_n578_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n933_), .A2(new_n205_), .A3(new_n577_), .A4(new_n913_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1353gat));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AND2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  NOR4_X1   g743(.A1(new_n934_), .A2(new_n639_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n934_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n640_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n947_), .B2(new_n943_), .ZN(G1354gat));
  XNOR2_X1  g747(.A(KEYINPUT127), .B(G218gat), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n934_), .A2(new_n688_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n946_), .A2(new_n526_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n949_), .ZN(G1355gat));
endmodule


