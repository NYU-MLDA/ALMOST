//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n206_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT22), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n218_), .B2(KEYINPUT78), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT22), .B(G169gat), .Z(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(KEYINPUT78), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT25), .B1(new_n207_), .B2(KEYINPUT74), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n223_), .B(new_n224_), .C1(new_n225_), .C2(KEYINPUT74), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(new_n216_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n204_), .A2(new_n227_), .A3(KEYINPUT24), .A4(new_n205_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n211_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n210_), .A2(KEYINPUT76), .A3(G183gat), .A4(G190gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n227_), .A2(KEYINPUT24), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n229_), .B1(new_n236_), .B2(KEYINPUT77), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n222_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(G15gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n244_), .B(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT80), .ZN(new_n250_));
  INV_X1    g049(.A(G134gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G127gat), .ZN(new_n252_));
  INV_X1    g051(.A(G127gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G134gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G120gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G113gat), .ZN(new_n257_));
  INV_X1    g056(.A(G113gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G120gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n255_), .A2(new_n260_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT79), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT31), .Z(new_n265_));
  OR2_X1    g064(.A1(new_n250_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n263_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n274_));
  NOR3_X1   g073(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT3), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n274_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n278_));
  INV_X1    g077(.A(G141gat), .ZN(new_n279_));
  INV_X1    g078(.A(G148gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(KEYINPUT3), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n270_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n280_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n284_), .A2(new_n271_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n268_), .A2(new_n287_), .A3(new_n269_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n267_), .B1(new_n290_), .B2(KEYINPUT94), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n281_), .A2(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n275_), .A2(new_n276_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n294_), .A2(new_n270_), .B1(new_n288_), .B2(new_n286_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT94), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n263_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT4), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT95), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n267_), .A2(new_n295_), .A3(KEYINPUT4), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n300_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G57gat), .B(G85gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT97), .ZN(new_n308_));
  INV_X1    g107(.A(G1gat), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n309_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n313_));
  INV_X1    g112(.A(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n306_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n304_), .A2(new_n305_), .A3(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n249_), .A2(KEYINPUT80), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n250_), .A2(new_n325_), .A3(new_n265_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n266_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n295_), .B2(new_n329_), .ZN(new_n330_));
  AND4_X1   g129(.A1(new_n328_), .A2(new_n283_), .A3(new_n329_), .A4(new_n289_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT82), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT28), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n295_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n332_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n333_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346_));
  AND2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT84), .B(KEYINPUT21), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n346_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(KEYINPUT21), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n345_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G197gat), .B(G204gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT84), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n354_), .A3(KEYINPUT85), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n356_), .B1(new_n361_), .B2(new_n344_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n343_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n344_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n352_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT85), .B1(new_n360_), .B2(new_n354_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n344_), .B1(new_n366_), .B2(new_n356_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(KEYINPUT86), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G233gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT83), .A2(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(KEYINPUT83), .A2(G228gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n295_), .B2(new_n329_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT87), .B1(new_n369_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n374_), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n363_), .A4(new_n368_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n353_), .A2(new_n362_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n375_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n342_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n342_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n340_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n389_), .B(new_n340_), .C1(new_n386_), .C2(KEYINPUT88), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n388_), .A2(new_n393_), .A3(new_n342_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n389_), .A2(new_n340_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n386_), .A2(KEYINPUT88), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n388_), .B2(new_n342_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n396_), .A2(KEYINPUT89), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n390_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT98), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n206_), .B1(new_n220_), .B2(G176gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT91), .ZN(new_n403_));
  INV_X1    g202(.A(new_n214_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n232_), .A2(new_n233_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n404_), .C1(new_n405_), .C2(new_n230_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT91), .B1(new_n234_), .B2(new_n214_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n402_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT25), .B(G183gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n223_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n412_), .A2(new_n235_), .A3(new_n213_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n383_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n237_), .A2(new_n239_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n222_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n363_), .A2(new_n368_), .ZN(new_n418_));
  OAI211_X1 g217(.A(KEYINPUT20), .B(new_n414_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n408_), .A2(new_n413_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n383_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n417_), .A2(new_n418_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n422_), .A3(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT93), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n424_), .A2(new_n430_), .A3(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(KEYINPUT27), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n419_), .A2(new_n423_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n422_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n240_), .A2(new_n369_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n408_), .A2(new_n383_), .A3(new_n413_), .ZN(new_n444_));
  NOR4_X1   g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n425_), .A4(new_n423_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n425_), .B1(new_n240_), .B2(new_n369_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n422_), .B1(new_n446_), .B2(new_n414_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n439_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n437_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT27), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n438_), .A2(new_n442_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n400_), .A2(new_n401_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n401_), .B1(new_n400_), .B2(new_n451_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n327_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n266_), .A2(new_n326_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n438_), .A2(new_n442_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n450_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n400_), .A2(new_n458_), .A3(new_n323_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n395_), .A2(new_n399_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n390_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n319_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n299_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n322_), .A2(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n304_), .A2(KEYINPUT33), .A3(new_n305_), .A4(new_n319_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n448_), .A3(new_n437_), .A4(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT32), .B(new_n436_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n424_), .A2(new_n430_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n323_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n460_), .A2(new_n461_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n455_), .B1(new_n459_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n454_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G29gat), .B(G36gat), .Z(new_n476_));
  XOR2_X1   g275(.A(G43gat), .B(G50gat), .Z(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n309_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G8gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n478_), .A2(new_n486_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT72), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n478_), .B(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n491_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n487_), .A2(new_n495_), .A3(new_n490_), .A4(new_n488_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G141gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .A4(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n504_), .B(KEYINPUT73), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n475_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n486_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n514_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n511_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G127gat), .B(G155gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT16), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(KEYINPUT71), .A2(KEYINPUT17), .ZN(new_n527_));
  OR3_X1    g326(.A1(new_n522_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  MUX2_X1   g327(.A(new_n527_), .B(KEYINPUT17), .S(new_n526_), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT64), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(KEYINPUT64), .A3(new_n533_), .ZN(new_n537_));
  AOI21_X1  g336(.A(G106gat), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT6), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT9), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G85gat), .B(G92gat), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n540_), .B(new_n542_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n538_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n544_), .B(KEYINPUT65), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT8), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n549_));
  OR3_X1    g348(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n540_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n546_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n480_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n478_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT70), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n555_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n564_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n563_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n568_), .B(KEYINPUT36), .Z(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT37), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT37), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n531_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT66), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n554_), .B2(new_n520_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n538_), .A2(new_n545_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n540_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT65), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n544_), .B(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT8), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n547_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n581_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(KEYINPUT66), .A3(new_n519_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n554_), .A2(new_n520_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n587_), .B2(new_n519_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n587_), .B2(new_n519_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n554_), .A2(KEYINPUT12), .A3(new_n520_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G120gat), .B(G148gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n592_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n578_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n509_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n613_), .A2(G1gat), .A3(new_n324_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n616_));
  INV_X1    g415(.A(new_n475_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n575_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n611_), .A2(new_n504_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n531_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n324_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n615_), .A2(new_n616_), .A3(new_n623_), .ZN(G1324gat));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n458_), .A3(new_n621_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n625_), .A2(G8gat), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n625_), .B2(G8gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n458_), .A2(new_n482_), .ZN(new_n629_));
  OAI22_X1  g428(.A1(new_n627_), .A2(new_n628_), .B1(new_n613_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n630_), .B(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n622_), .B2(new_n455_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n455_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n246_), .ZN(new_n639_));
  OAI22_X1  g438(.A1(new_n636_), .A2(new_n637_), .B1(new_n613_), .B2(new_n639_), .ZN(G1326gat));
  OR3_X1    g439(.A1(new_n613_), .A2(G22gat), .A3(new_n400_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n622_), .B2(new_n400_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT103), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n644_), .B(G22gat), .C1(new_n622_), .C2(new_n400_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n646_));
  AND3_X1   g445(.A1(new_n643_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n641_), .B1(new_n647_), .B2(new_n648_), .ZN(G1327gat));
  NAND2_X1  g448(.A1(new_n618_), .A2(new_n531_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT104), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n610_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n509_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n323_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n531_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n620_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n576_), .A2(new_n577_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n475_), .B2(new_n660_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT43), .B(new_n659_), .C1(new_n454_), .C2(new_n474_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT44), .B(new_n657_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n324_), .A2(new_n314_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n655_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n458_), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n451_), .A2(G36gat), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n509_), .A2(new_n672_), .A3(new_n652_), .A4(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n507_), .A2(new_n508_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT99), .B1(new_n475_), .B2(new_n506_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n652_), .B(new_n673_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT45), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n674_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n671_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  OAI21_X1  g483(.A(new_n242_), .B1(new_n653_), .B2(new_n455_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n665_), .A2(G43gat), .A3(new_n638_), .A4(new_n666_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1330gat));
  INV_X1    g489(.A(new_n400_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G50gat), .B1(new_n654_), .B2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(G50gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n667_), .B2(new_n693_), .ZN(G1331gat));
  INV_X1    g493(.A(new_n504_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n610_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n617_), .A2(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n697_), .A2(KEYINPUT106), .A3(new_n578_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT106), .B1(new_n697_), .B2(new_n578_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n323_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  AND4_X1   g504(.A1(new_n505_), .A2(new_n619_), .A3(new_n610_), .A4(new_n656_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n324_), .A2(new_n705_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n704_), .A2(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(G1332gat));
  NOR2_X1   g507(.A1(new_n451_), .A2(G64gat), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT108), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n700_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n458_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G64gat), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(KEYINPUT48), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(KEYINPUT48), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n700_), .A2(new_n717_), .A3(new_n638_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n706_), .A2(new_n638_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G71gat), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT49), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT49), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1334gat));
  NOR2_X1   g522(.A1(new_n400_), .A2(G78gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT109), .Z(new_n725_));
  NAND2_X1  g524(.A1(new_n700_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n706_), .A2(new_n691_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G78gat), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT50), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT50), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n617_), .A2(new_n651_), .A3(new_n696_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n323_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n661_), .A2(new_n662_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n611_), .A2(new_n504_), .A3(new_n656_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n323_), .A2(G85gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT111), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n737_), .B1(new_n740_), .B2(new_n742_), .ZN(G1336gat));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n736_), .A2(new_n744_), .A3(new_n458_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n740_), .A2(new_n458_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(new_n746_), .ZN(G1337gat));
  AND2_X1   g546(.A1(new_n536_), .A2(new_n537_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n638_), .B(new_n749_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n738_), .A2(new_n638_), .A3(new_n739_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G99gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(G1338gat));
  INV_X1    g554(.A(G106gat), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n691_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n691_), .B(new_n739_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n760_));
  AND4_X1   g559(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .A4(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n760_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n756_), .B1(new_n762_), .B2(KEYINPUT114), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n759_), .A2(new_n763_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n757_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n757_), .B(new_n767_), .C1(new_n761_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  NAND3_X1  g568(.A1(new_n578_), .A2(new_n505_), .A3(new_n611_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n500_), .B1(new_n493_), .B2(new_n490_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n503_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n606_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT117), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n606_), .A2(new_n779_), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n597_), .A2(KEYINPUT55), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .A4(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n580_), .A2(new_n594_), .A3(new_n596_), .A4(new_n588_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n782_), .A2(new_n784_), .B1(new_n591_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n602_), .B1(new_n786_), .B2(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n591_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n792_), .A3(KEYINPUT56), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n792_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT116), .B(KEYINPUT56), .C1(new_n787_), .C2(new_n792_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n695_), .A2(new_n604_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n781_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n773_), .B1(new_n801_), .B2(new_n618_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n618_), .A2(new_n773_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n800_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n602_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n796_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n795_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n807_), .B1(new_n814_), .B2(new_n793_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT119), .B(new_n804_), .C1(new_n815_), .C2(new_n781_), .ZN(new_n816_));
  OR3_X1    g615(.A1(new_n795_), .A2(KEYINPUT118), .A3(new_n796_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(KEYINPUT118), .A3(new_n793_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n776_), .A2(new_n603_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n659_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n817_), .A2(new_n818_), .A3(KEYINPUT58), .A4(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n802_), .A2(new_n806_), .A3(new_n816_), .A4(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n772_), .B1(new_n825_), .B2(new_n531_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n323_), .B(new_n638_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n826_), .A2(KEYINPUT120), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT120), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n258_), .A4(new_n504_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n825_), .A2(new_n531_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n772_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n827_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT59), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n505_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n258_), .ZN(G1340gat));
  XOR2_X1   g638(.A(KEYINPUT121), .B(G120gat), .Z(new_n840_));
  OR2_X1    g639(.A1(new_n840_), .A2(KEYINPUT60), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n611_), .B2(KEYINPUT60), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n828_), .A2(new_n829_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n611_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n840_), .ZN(G1341gat));
  NAND4_X1  g644(.A1(new_n828_), .A2(new_n829_), .A3(new_n253_), .A4(new_n656_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n531_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n253_), .ZN(G1342gat));
  NAND4_X1  g647(.A1(new_n828_), .A2(new_n829_), .A3(new_n251_), .A4(new_n618_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n659_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n251_), .ZN(G1343gat));
  NOR4_X1   g650(.A1(new_n638_), .A2(new_n400_), .A3(new_n458_), .A4(new_n324_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n504_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n610_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n854_), .B2(new_n656_), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n826_), .A2(KEYINPUT122), .A3(new_n531_), .A4(new_n853_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n806_), .A2(new_n816_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n575_), .B1(new_n815_), .B2(new_n781_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n866_), .A2(new_n773_), .B1(new_n823_), .B2(new_n822_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n656_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n656_), .B(new_n852_), .C1(new_n868_), .C2(new_n772_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT122), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n854_), .A2(new_n861_), .A3(new_n656_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n859_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(new_n872_), .ZN(G1346gat));
  INV_X1    g672(.A(new_n854_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G162gat), .B1(new_n874_), .B2(new_n659_), .ZN(new_n875_));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n854_), .A2(new_n876_), .A3(new_n618_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n451_), .A2(new_n323_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n638_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n695_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n400_), .B1(new_n882_), .B2(KEYINPUT123), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(KEYINPUT123), .B2(new_n882_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n217_), .B1(new_n833_), .B2(new_n884_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(KEYINPUT125), .A3(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n826_), .A2(new_n691_), .A3(new_n880_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n695_), .A2(new_n220_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n886_), .B(KEYINPUT125), .Z(new_n892_));
  OAI211_X1 g691(.A(new_n888_), .B(new_n891_), .C1(new_n885_), .C2(new_n892_), .ZN(G1348gat));
  NAND4_X1  g692(.A1(new_n833_), .A2(new_n400_), .A3(new_n638_), .A4(new_n879_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n894_), .A2(new_n216_), .A3(new_n611_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G176gat), .B1(new_n889_), .B2(new_n610_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1349gat));
  NOR3_X1   g696(.A1(new_n894_), .A2(new_n409_), .A3(new_n531_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G183gat), .B1(new_n889_), .B2(new_n656_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n894_), .B2(new_n659_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n223_), .A3(new_n618_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  NAND3_X1  g702(.A1(new_n455_), .A2(new_n879_), .A3(new_n691_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n504_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n610_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g708(.A(new_n531_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT126), .Z(new_n913_));
  XNOR2_X1  g712(.A(new_n911_), .B(new_n913_), .ZN(G1354gat));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n905_), .B2(new_n660_), .ZN(new_n917_));
  NOR4_X1   g716(.A1(new_n826_), .A2(G218gat), .A3(new_n575_), .A4(new_n904_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n905_), .A2(new_n916_), .A3(new_n618_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n826_), .A2(new_n659_), .A3(new_n904_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n920_), .B(KEYINPUT127), .C1(new_n921_), .C2(new_n916_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n922_), .ZN(G1355gat));
endmodule


