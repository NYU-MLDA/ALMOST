//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n212_), .A2(KEYINPUT9), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n208_), .B1(KEYINPUT9), .B2(new_n202_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT65), .ZN(new_n223_));
  XOR2_X1   g022(.A(G71gat), .B(G78gat), .Z(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(KEYINPUT11), .B2(new_n221_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n223_), .B(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n220_), .B(new_n226_), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT12), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT12), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G230gat), .A2(G233gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n227_), .A2(new_n232_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G120gat), .B(G148gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT5), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G176gat), .B(G204gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT13), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(KEYINPUT13), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G29gat), .B(G36gat), .Z(new_n247_));
  XOR2_X1   g046(.A(G43gat), .B(G50gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT15), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n220_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT34), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT66), .B(KEYINPUT35), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n249_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n220_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n254_), .A2(new_n255_), .ZN(new_n259_));
  OR3_X1    g058(.A1(new_n251_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G190gat), .B(G218gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT67), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G134gat), .B(G162gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT36), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT68), .Z(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT69), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n260_), .A2(new_n271_), .A3(new_n261_), .A4(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(KEYINPUT70), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT70), .B1(new_n270_), .B2(new_n272_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n265_), .B(KEYINPUT36), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n274_), .A2(new_n275_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT37), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT71), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n275_), .A2(new_n278_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n282_), .B(KEYINPUT37), .C1(new_n283_), .C2(new_n274_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n278_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n280_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT72), .B(G15gat), .ZN(new_n289_));
  INV_X1    g088(.A(G22gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT73), .B(G1gat), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G8gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(KEYINPUT14), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT74), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(new_n226_), .Z(new_n300_));
  INV_X1    g099(.A(KEYINPUT17), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G155gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G183gat), .B(G211gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  OR3_X1    g105(.A1(new_n300_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(KEYINPUT17), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n288_), .A2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n311_), .A2(KEYINPUT76), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(KEYINPUT76), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n246_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n295_), .B(new_n296_), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n249_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n297_), .A2(new_n257_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n297_), .A2(KEYINPUT77), .A3(new_n257_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n297_), .A2(new_n250_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n324_), .A3(new_n320_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G141gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G169gat), .B(G197gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OR3_X1    g131(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  INV_X1    g139(.A(G155gat), .ZN(new_n341_));
  INV_X1    g140(.A(G162gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n343_), .A2(new_n344_), .B1(G155gat), .B2(G162gat), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n334_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(new_n344_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT29), .B1(new_n346_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(G218gat), .ZN(new_n358_));
  INV_X1    g157(.A(G218gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(G211gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT86), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(G211gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(G218gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G197gat), .B(G204gat), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n361_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n361_), .A2(new_n365_), .B1(KEYINPUT85), .B2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT21), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(KEYINPUT85), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n364_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT21), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n356_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n369_), .A2(new_n377_), .A3(new_n375_), .ZN(new_n378_));
  INV_X1    g177(.A(G228gat), .ZN(new_n379_));
  INV_X1    g178(.A(G233gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(new_n378_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n361_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n374_), .B1(new_n373_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n361_), .A2(new_n365_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT21), .B1(new_n386_), .B2(new_n370_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n388_), .B(new_n356_), .C1(new_n377_), .C2(new_n381_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n383_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n353_), .A2(new_n354_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n350_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n339_), .A2(new_n345_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT28), .B1(new_n400_), .B2(KEYINPUT29), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n398_), .A2(new_n402_), .A3(new_n399_), .A4(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G22gat), .B(G50gat), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n401_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n395_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n394_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n413_), .B(new_n391_), .C1(new_n383_), .C2(new_n389_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT87), .B1(new_n390_), .B2(new_n392_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n390_), .A2(KEYINPUT87), .A3(new_n392_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n394_), .A3(new_n408_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n420_), .A2(KEYINPUT88), .A3(new_n416_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n410_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G127gat), .B(G134gat), .Z(new_n426_));
  XOR2_X1   g225(.A(G113gat), .B(G120gat), .Z(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n400_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n426_), .B(new_n427_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(KEYINPUT4), .A3(new_n431_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(KEYINPUT4), .B2(new_n429_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n432_), .B1(new_n434_), .B2(new_n425_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G85gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT0), .B(G57gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n441_));
  INV_X1    g240(.A(new_n439_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n429_), .A2(KEYINPUT4), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n424_), .B1(new_n443_), .B2(new_n433_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n444_), .B2(new_n432_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n435_), .A2(KEYINPUT98), .A3(new_n439_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(KEYINPUT23), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT23), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(KEYINPUT80), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(G183gat), .A3(G190gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n458_), .A3(KEYINPUT23), .ZN(new_n459_));
  INV_X1    g258(.A(G183gat), .ZN(new_n460_));
  INV_X1    g259(.A(G190gat), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n455_), .A2(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n463_));
  INV_X1    g262(.A(G169gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G169gat), .A2(G176gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT25), .B1(new_n460_), .B2(KEYINPUT78), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(G183gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT26), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(new_n474_), .A3(new_n476_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n453_), .B1(G183gat), .B2(G190gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n456_), .A2(new_n458_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(new_n453_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n462_), .A2(new_n465_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G43gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(new_n428_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(G15gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT30), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT31), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n449_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G8gat), .B(G36gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT19), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(KEYINPUT20), .C1(new_n388_), .C2(new_n484_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT25), .B(G183gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G190gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n477_), .A2(G190gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n461_), .A2(KEYINPUT26), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT90), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n509_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n455_), .A2(new_n459_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n470_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n469_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n519_), .A2(KEYINPUT91), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(KEYINPUT91), .ZN(new_n521_));
  INV_X1    g320(.A(G176gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT22), .B(G169gat), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n520_), .A2(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G183gat), .A2(G190gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n524_), .B1(new_n483_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n388_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n508_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n462_), .A2(new_n465_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n480_), .A2(new_n483_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n530_), .B(new_n531_), .C1(new_n385_), .C2(new_n387_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n507_), .B1(new_n532_), .B2(KEYINPUT20), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n504_), .B(new_n506_), .C1(new_n529_), .C2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n518_), .B(new_n526_), .C1(new_n385_), .C2(new_n387_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n369_), .A2(new_n484_), .A3(new_n375_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n506_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT20), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT92), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n484_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT89), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n528_), .A3(new_n508_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n544_), .B2(new_n506_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n503_), .B1(new_n535_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n508_), .A2(new_n528_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n548_), .B2(new_n543_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n502_), .B(new_n534_), .C1(new_n549_), .C2(new_n540_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT27), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n535_), .A2(new_n545_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(KEYINPUT94), .A3(new_n502_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT100), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT100), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n551_), .A2(new_n557_), .A3(new_n554_), .A4(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT20), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n506_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n544_), .B2(new_n506_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n502_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n546_), .A2(KEYINPUT27), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT101), .B1(new_n559_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT101), .ZN(new_n566_));
  INV_X1    g365(.A(new_n564_), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n566_), .B(new_n567_), .C1(new_n556_), .C2(new_n558_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n423_), .B(new_n497_), .C1(new_n565_), .C2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n496_), .B(KEYINPUT82), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT95), .B1(new_n435_), .B2(new_n439_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT33), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n445_), .A2(KEYINPUT95), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n429_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n439_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT96), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT96), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n577_), .B(new_n578_), .C1(new_n425_), .C2(new_n434_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n503_), .A2(KEYINPUT32), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT97), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n553_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n562_), .A2(new_n582_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n446_), .A2(new_n585_), .A3(new_n447_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n423_), .B1(new_n581_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT99), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n423_), .B(new_n590_), .C1(new_n581_), .C2(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n422_), .A2(new_n448_), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n567_), .B(new_n593_), .C1(new_n556_), .C2(new_n558_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n570_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n332_), .B1(new_n569_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n314_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n292_), .B1(KEYINPUT102), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n449_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(KEYINPUT102), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n246_), .A2(new_n310_), .A3(new_n332_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n569_), .A2(new_n595_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n285_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n604_), .A2(KEYINPUT103), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT103), .B1(new_n604_), .B2(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n448_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(new_n565_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n568_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(G8gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n314_), .A2(new_n596_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT104), .ZN(new_n616_));
  OAI21_X1  g415(.A(G8gat), .B1(new_n608_), .B2(new_n613_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n621_), .B(new_n623_), .ZN(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n608_), .B2(new_n570_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  INV_X1    g425(.A(new_n570_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n597_), .A2(new_n490_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1326gat));
  NAND3_X1  g428(.A1(new_n597_), .A2(new_n290_), .A3(new_n422_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G22gat), .B1(new_n608_), .B2(new_n423_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(G1327gat));
  NAND2_X1  g434(.A1(new_n310_), .A2(new_n285_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n246_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n596_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(G29gat), .B1(new_n639_), .B2(new_n449_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n310_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(new_n246_), .A3(new_n332_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n604_), .B2(new_n288_), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT43), .B(new_n287_), .C1(new_n569_), .C2(new_n595_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT44), .B(new_n642_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n449_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n640_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n613_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n613_), .A2(new_n653_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n658_), .A2(new_n659_), .A3(new_n639_), .A4(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n663_), .B2(new_n638_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n613_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n648_), .A2(new_n666_), .A3(new_n649_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(new_n667_), .B2(G36gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT110), .B1(new_n668_), .B2(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT109), .B(new_n665_), .C1(new_n667_), .C2(G36gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n667_), .A2(G36gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n665_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT109), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n668_), .A2(new_n671_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n678_), .A2(KEYINPUT110), .A3(new_n670_), .A4(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n674_), .A2(new_n680_), .ZN(G1329gat));
  INV_X1    g480(.A(new_n496_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n650_), .A2(G43gat), .A3(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT111), .B(G43gat), .Z(new_n684_));
  OAI21_X1  g483(.A(new_n684_), .B1(new_n638_), .B2(new_n570_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n639_), .B2(new_n422_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n422_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n650_), .B2(new_n689_), .ZN(G1331gat));
  INV_X1    g489(.A(new_n246_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n332_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n569_), .B2(new_n595_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n449_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n606_), .A2(new_n607_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n691_), .A2(new_n693_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n641_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n448_), .A2(KEYINPUT112), .ZN(new_n701_));
  MUX2_X1   g500(.A(KEYINPUT112), .B(new_n701_), .S(G57gat), .Z(new_n702_));
  AOI21_X1  g501(.A(new_n696_), .B1(new_n700_), .B2(new_n702_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n695_), .A2(new_n704_), .A3(new_n658_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n700_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G64gat), .B1(new_n706_), .B2(new_n657_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT48), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT48), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n700_), .B2(new_n627_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT49), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n695_), .A2(new_n711_), .A3(new_n627_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n695_), .A2(new_n716_), .A3(new_n422_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n700_), .A2(new_n422_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G78gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT50), .B(new_n716_), .C1(new_n700_), .C2(new_n422_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT113), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n636_), .A2(new_n691_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n694_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n449_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n310_), .B(new_n698_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT114), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n448_), .A2(new_n212_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n213_), .A3(new_n666_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n658_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n213_), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n728_), .B2(new_n570_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n216_), .A3(new_n682_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g537(.A(G106gat), .B1(new_n728_), .B2(new_n423_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT52), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n726_), .A2(new_n217_), .A3(new_n422_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g542(.A(KEYINPUT120), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n666_), .A2(new_n422_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n448_), .A2(new_n496_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT59), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n240_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n232_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n228_), .A2(new_n752_), .A3(new_n230_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(KEYINPUT55), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT115), .B1(new_n233_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n754_), .A2(new_n758_), .A3(KEYINPUT55), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n238_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n238_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n751_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n320_), .B1(new_n315_), .B2(new_n249_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n328_), .B1(new_n767_), .B2(new_n324_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n330_), .B(new_n243_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n605_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(KEYINPUT117), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n760_), .A2(new_n774_), .A3(KEYINPUT56), .A4(new_n238_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n763_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n766_), .A2(new_n768_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n329_), .A2(new_n240_), .A3(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT116), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n287_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n779_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n782_), .A2(new_n783_), .B1(new_n771_), .B2(new_n770_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n772_), .B1(new_n784_), .B2(KEYINPUT119), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n783_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n770_), .A2(new_n771_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(KEYINPUT119), .A3(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n310_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n691_), .A2(new_n641_), .A3(new_n287_), .A4(new_n332_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n750_), .B1(new_n789_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n786_), .A2(new_n772_), .A3(new_n787_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n310_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n793_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n749_), .B1(new_n797_), .B2(new_n748_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n744_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n792_), .B1(new_n795_), .B2(new_n310_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT59), .B1(new_n800_), .B2(new_n747_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n780_), .A2(new_n781_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(new_n288_), .A3(new_n783_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n787_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n802_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n784_), .A2(KEYINPUT119), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n772_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n792_), .B1(new_n808_), .B2(new_n310_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT120), .B(new_n801_), .C1(new_n809_), .C2(new_n750_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n799_), .A2(G113gat), .A3(new_n810_), .A4(new_n693_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n800_), .A2(new_n747_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n693_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT118), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n811_), .A2(new_n814_), .ZN(G1340gat));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n691_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n812_), .B(new_n817_), .C1(KEYINPUT60), .C2(new_n816_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n794_), .A2(new_n798_), .A3(new_n691_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n816_), .ZN(G1341gat));
  NAND3_X1  g619(.A1(new_n799_), .A2(new_n641_), .A3(new_n810_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G127gat), .ZN(new_n822_));
  INV_X1    g621(.A(G127gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n812_), .A2(new_n823_), .A3(new_n641_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1342gat));
  NAND4_X1  g624(.A1(new_n799_), .A2(G134gat), .A3(new_n810_), .A4(new_n288_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G134gat), .B1(new_n812_), .B2(new_n285_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT121), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1343gat));
  NOR2_X1   g628(.A1(new_n800_), .A2(new_n627_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n830_), .A2(new_n449_), .A3(new_n422_), .A4(new_n657_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n332_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(new_n347_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n691_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n348_), .ZN(G1345gat));
  NOR2_X1   g634(.A1(new_n831_), .A2(new_n310_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT61), .B(G155gat), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n836_), .B(new_n837_), .Z(G1346gat));
  OAI21_X1  g637(.A(G162gat), .B1(new_n831_), .B2(new_n287_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n285_), .A2(new_n342_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n831_), .B2(new_n840_), .ZN(G1347gat));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n789_), .A2(new_n793_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n657_), .A2(new_n449_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n570_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n423_), .A3(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n332_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n842_), .B1(new_n848_), .B2(new_n464_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n523_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT62), .B(G169gat), .C1(new_n847_), .C2(new_n332_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(G1348gat));
  NOR2_X1   g651(.A1(new_n800_), .A2(new_n422_), .ZN(new_n853_));
  AND4_X1   g652(.A1(G176gat), .A2(new_n853_), .A3(new_n246_), .A4(new_n846_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n809_), .A2(new_n422_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n246_), .A3(new_n846_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n522_), .ZN(G1349gat));
  NOR4_X1   g656(.A1(new_n845_), .A2(new_n570_), .A3(new_n509_), .A4(new_n310_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n853_), .A2(new_n641_), .A3(new_n846_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n855_), .A2(new_n858_), .B1(new_n859_), .B2(new_n460_), .ZN(G1350gat));
  NAND4_X1  g659(.A1(new_n843_), .A2(new_n423_), .A3(new_n288_), .A4(new_n846_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n861_), .A2(new_n862_), .A3(G190gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n861_), .B2(G190gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n285_), .B1(new_n515_), .B2(new_n512_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT123), .Z(new_n866_));
  OAI22_X1  g665(.A1(new_n863_), .A2(new_n864_), .B1(new_n847_), .B2(new_n866_), .ZN(G1351gat));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n800_), .A2(new_n845_), .A3(new_n627_), .A4(new_n423_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n693_), .ZN(new_n870_));
  INV_X1    g669(.A(G197gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n868_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n871_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n869_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n693_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(G1352gat));
  NAND2_X1  g674(.A1(new_n869_), .A2(new_n246_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g676(.A1(new_n830_), .A2(new_n422_), .A3(new_n844_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n310_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT125), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n869_), .A2(new_n882_), .A3(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n881_), .A2(new_n885_), .A3(new_n883_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1354gat));
  OAI21_X1  g688(.A(new_n359_), .B1(new_n878_), .B2(new_n605_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n287_), .A2(new_n359_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT126), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n869_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n890_), .A2(KEYINPUT127), .A3(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1355gat));
endmodule


