//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT72), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  INV_X1    g005(.A(G43gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G50gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n206_), .B(G43gat), .ZN(new_n210_));
  INV_X1    g009(.A(G50gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT15), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G85gat), .B(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT66), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT66), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n217_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n219_), .A2(new_n221_), .ZN(new_n231_));
  AOI211_X1 g030(.A(new_n230_), .B(new_n215_), .C1(new_n228_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n220_), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n225_), .B(new_n236_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n215_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n232_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n229_), .B1(new_n242_), .B2(KEYINPUT8), .ZN(new_n243_));
  OR2_X1    g042(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n244_), .A2(G85gat), .A3(G92gat), .A4(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n215_), .B2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n234_), .A2(KEYINPUT10), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT10), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G99gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(G106gat), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  NOR4_X1   g050(.A1(new_n247_), .A2(new_n222_), .A3(new_n223_), .A4(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT68), .B1(new_n243_), .B2(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n219_), .A2(new_n221_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n236_), .A2(new_n225_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n240_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n230_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n239_), .A2(KEYINPUT67), .A3(new_n240_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT8), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n224_), .A2(new_n228_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n216_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n252_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n214_), .B1(new_n253_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n205_), .B1(new_n265_), .B2(KEYINPUT73), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT15), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n213_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n259_), .A2(new_n261_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n252_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n263_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AOI211_X1 g070(.A(KEYINPUT68), .B(new_n252_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n274_));
  INV_X1    g073(.A(new_n213_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n262_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n266_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n253_), .A2(new_n264_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n268_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n281_), .A2(new_n283_), .A3(new_n205_), .A4(new_n274_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G134gat), .ZN(new_n286_));
  INV_X1    g085(.A(G162gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT36), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n278_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT36), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n291_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT37), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n278_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n205_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n273_), .B2(new_n282_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(new_n277_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n302_), .B2(new_n294_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G8gat), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT75), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G1gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n306_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n307_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n306_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G8gat), .A3(new_n314_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G231gat), .ZN(new_n321_));
  INV_X1    g120(.A(G233gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G57gat), .B(G64gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT11), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G71gat), .B(G78gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n325_), .A2(KEYINPUT11), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n323_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n324_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n324_), .B2(new_n331_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G155gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G183gat), .B(G211gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n340_), .A2(KEYINPUT17), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n334_), .A2(KEYINPUT77), .A3(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n340_), .A2(KEYINPUT17), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n334_), .A2(new_n341_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n305_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n351_));
  INV_X1    g150(.A(new_n330_), .ZN(new_n352_));
  OAI211_X1 g151(.A(KEYINPUT12), .B(new_n352_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n352_), .B1(new_n243_), .B2(new_n252_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT69), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT69), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n262_), .A2(new_n330_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G230gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT64), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n359_), .A2(KEYINPUT70), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT70), .B1(new_n359_), .B2(new_n362_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n353_), .B(new_n358_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n354_), .A2(new_n359_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n361_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G120gat), .B(G148gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT5), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G176gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G204gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n365_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n365_), .A2(new_n367_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n371_), .B(KEYINPUT71), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n351_), .B(new_n372_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n365_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT13), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n213_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n317_), .A2(new_n319_), .A3(new_n213_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G229gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(G8gat), .B1(new_n318_), .B2(new_n314_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n315_), .A2(new_n306_), .A3(new_n316_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n381_), .B1(new_n268_), .B2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n385_), .B(KEYINPUT79), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n384_), .A2(KEYINPUT78), .A3(new_n386_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G113gat), .B(G141gat), .ZN(new_n398_));
  INV_X1    g197(.A(G169gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(G197gat), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n389_), .A2(new_n396_), .A3(new_n397_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT80), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT78), .B1(new_n384_), .B2(new_n386_), .ZN(new_n405_));
  AOI211_X1 g204(.A(new_n388_), .B(new_n385_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n396_), .A4(new_n402_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n396_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n401_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n380_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n419_));
  OR2_X1    g218(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n418_), .A2(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT24), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n416_), .B1(new_n422_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT23), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n425_), .A2(new_n426_), .ZN(new_n437_));
  AND2_X1   g236(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n438_));
  AND2_X1   g237(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n440_));
  OAI22_X1  g239(.A1(new_n417_), .A2(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G176gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n399_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT24), .A3(new_n423_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(KEYINPUT87), .A3(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n428_), .A2(new_n436_), .A3(new_n437_), .A4(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G211gat), .B(G218gat), .ZN(new_n447_));
  INV_X1    g246(.A(G204gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT85), .B1(new_n448_), .B2(G197gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(KEYINPUT21), .A3(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G197gat), .B(G204gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n447_), .A2(KEYINPUT21), .ZN(new_n453_));
  XOR2_X1   g252(.A(G197gat), .B(G204gat), .Z(new_n454_));
  NAND4_X1  g253(.A1(new_n454_), .A2(KEYINPUT21), .A3(new_n447_), .A4(new_n449_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n431_), .A2(new_n434_), .A3(new_n432_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n429_), .A2(KEYINPUT23), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G183gat), .ZN(new_n460_));
  INV_X1    g259(.A(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465_));
  NAND2_X1  g264(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n442_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n469_), .A3(new_n423_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n446_), .A2(new_n456_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT19), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(KEYINPUT20), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n456_), .A2(KEYINPUT86), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n452_), .A2(new_n455_), .A3(new_n477_), .A4(new_n453_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n441_), .A2(new_n444_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT81), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT81), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n441_), .A2(new_n481_), .A3(new_n444_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n480_), .A2(new_n482_), .A3(new_n437_), .A4(new_n459_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n436_), .A2(new_n462_), .ZN(new_n484_));
  AOI21_X1  g283(.A(G176gat), .B1(KEYINPUT83), .B2(KEYINPUT22), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G169gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n476_), .A2(new_n478_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n475_), .A2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n436_), .A2(new_n445_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n479_), .A2(new_n416_), .B1(new_n426_), .B2(new_n425_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n424_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n490_), .A2(new_n491_), .B1(new_n492_), .B2(new_n469_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n493_), .B2(new_n456_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n476_), .A2(new_n483_), .A3(new_n487_), .A4(new_n478_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n446_), .A2(new_n470_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497_));
  INV_X1    g296(.A(new_n456_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n494_), .A2(KEYINPUT20), .A3(new_n495_), .A4(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n489_), .B1(new_n500_), .B2(new_n473_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT18), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G64gat), .ZN(new_n504_));
  INV_X1    g303(.A(G92gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT90), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508_));
  INV_X1    g307(.A(new_n506_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n497_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n510_));
  AOI211_X1 g309(.A(KEYINPUT89), .B(new_n456_), .C1(new_n446_), .C2(new_n470_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n495_), .A2(KEYINPUT20), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n474_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n508_), .B(new_n509_), .C1(new_n514_), .C2(new_n489_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n501_), .A2(new_n506_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT96), .B(KEYINPUT27), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G134gat), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G120gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G113gat), .ZN(new_n523_));
  INV_X1    g322(.A(G113gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G120gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n521_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(new_n525_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT84), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT3), .ZN(new_n535_));
  INV_X1    g334(.A(G141gat), .ZN(new_n536_));
  INV_X1    g335(.A(G148gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G141gat), .A2(G148gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT2), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(G155gat), .A2(G162gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G155gat), .A2(G162gat), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(KEYINPUT1), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT1), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(G155gat), .A3(G162gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n551_), .A3(new_n545_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G141gat), .B(G148gat), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n554_), .A3(KEYINPUT91), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n534_), .A2(new_n555_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n544_), .A2(new_n547_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n557_), .A2(new_n530_), .A3(KEYINPUT91), .A4(new_n533_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n558_), .A3(KEYINPUT4), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G225gat), .A2(G233gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(KEYINPUT4), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n561_), .B2(new_n534_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n556_), .A2(new_n558_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n560_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n559_), .A2(KEYINPUT92), .A3(new_n562_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G1gat), .B(G29gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G85gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n565_), .A2(new_n574_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(G228gat), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n322_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT29), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n557_), .A2(new_n581_), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n580_), .B(new_n582_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n456_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G78gat), .B(G106gat), .ZN(new_n586_));
  INV_X1    g385(.A(G22gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n583_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n476_), .A2(new_n478_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n580_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n582_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n590_), .B1(new_n594_), .B2(new_n584_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n548_), .A2(new_n554_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT28), .B1(new_n596_), .B2(KEYINPUT29), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT28), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n557_), .A2(new_n598_), .A3(new_n581_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n597_), .A2(new_n211_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n211_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n589_), .A2(new_n595_), .A3(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n600_), .A2(new_n601_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n588_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n594_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G15gat), .B(G43gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT31), .ZN(new_n609_));
  INV_X1    g408(.A(new_n534_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G71gat), .B(G99gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT30), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G227gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n483_), .A2(new_n487_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n534_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n609_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n611_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n618_), .B1(new_n614_), .B2(new_n622_), .ZN(new_n625_));
  OAI22_X1  g424(.A1(new_n603_), .A2(new_n607_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n602_), .B1(new_n589_), .B2(new_n595_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n614_), .A2(new_n622_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n618_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n605_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n627_), .A2(new_n630_), .A3(new_n623_), .A4(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n578_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(KEYINPUT95), .A2(KEYINPUT20), .ZN(new_n634_));
  NAND2_X1  g433(.A1(KEYINPUT95), .A2(KEYINPUT20), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n471_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n473_), .B1(new_n636_), .B2(new_n488_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n500_), .B2(new_n473_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n509_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n516_), .A3(KEYINPUT27), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n519_), .A2(new_n633_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n506_), .A2(KEYINPUT32), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n501_), .A2(new_n642_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n578_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n507_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n561_), .A2(new_n534_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n559_), .A2(new_n560_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n566_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n649_), .B(new_n575_), .C1(new_n650_), .C2(new_n560_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n577_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n577_), .A2(new_n652_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n577_), .A2(KEYINPUT94), .A3(new_n652_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n646_), .B1(new_n647_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n624_), .A2(new_n625_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n603_), .A2(new_n607_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n641_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n350_), .A2(new_n415_), .A3(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT97), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n578_), .A3(new_n311_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT38), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n379_), .A2(KEYINPUT98), .A3(new_n413_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT98), .B1(new_n379_), .B2(new_n413_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n349_), .A2(new_n303_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n664_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n578_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT99), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n668_), .A2(new_n676_), .ZN(G1324gat));
  NAND2_X1  g476(.A1(new_n519_), .A2(new_n640_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n666_), .A2(new_n306_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G8gat), .B1(new_n673_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT39), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n673_), .B2(new_n661_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT41), .Z(new_n686_));
  INV_X1    g485(.A(G15gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n666_), .A2(new_n687_), .A3(new_n660_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1326gat));
  INV_X1    g488(.A(new_n662_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n666_), .A2(new_n587_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G22gat), .B1(new_n673_), .B2(new_n662_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT42), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n349_), .A2(new_n303_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT100), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n415_), .A4(new_n664_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n695_), .A2(KEYINPUT100), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n349_), .B2(new_n303_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n415_), .B(new_n664_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT101), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n578_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n334_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n345_), .B2(new_n342_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n669_), .A2(new_n670_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT74), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n278_), .A2(new_n284_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n293_), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n711_), .B(new_n297_), .C1(new_n713_), .C2(new_n299_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT37), .B1(new_n303_), .B2(KEYINPUT74), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n664_), .B(new_n710_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n710_), .B1(new_n305_), .B2(new_n664_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n709_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT44), .B(new_n709_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n578_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n706_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  NAND3_X1  g525(.A1(new_n721_), .A2(new_n678_), .A3(new_n722_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n721_), .A2(KEYINPUT102), .A3(new_n678_), .A4(new_n722_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(G36gat), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n698_), .A2(new_n703_), .A3(new_n732_), .A4(new_n678_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(KEYINPUT46), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n731_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT104), .B(KEYINPUT46), .Z(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n736_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  NOR4_X1   g542(.A1(new_n738_), .A2(new_n739_), .A3(KEYINPUT105), .A4(new_n741_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n735_), .B1(new_n743_), .B2(new_n744_), .ZN(G1329gat));
  NAND2_X1  g544(.A1(KEYINPUT106), .A2(G43gat), .ZN(new_n746_));
  OR2_X1    g545(.A1(KEYINPUT106), .A2(G43gat), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n747_), .C1(new_n704_), .C2(new_n661_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n660_), .A2(G43gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n723_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g550(.A(G50gat), .B1(new_n723_), .B2(new_n662_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n705_), .A2(new_n211_), .A3(new_n690_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n379_), .A2(new_n413_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n664_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n672_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT107), .Z(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT108), .B(G57gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n578_), .A3(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT109), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n350_), .A2(new_n756_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n578_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1332gat));
  INV_X1    g563(.A(G64gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n758_), .B2(new_n678_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT48), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n765_), .A3(new_n678_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1333gat));
  INV_X1    g568(.A(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n758_), .B2(new_n660_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT49), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n762_), .A2(new_n770_), .A3(new_n660_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1334gat));
  INV_X1    g573(.A(G78gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n758_), .B2(new_n690_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT50), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n762_), .A2(new_n775_), .A3(new_n690_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1335gat));
  NAND2_X1  g578(.A1(new_n696_), .A2(new_n756_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n578_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n349_), .B(new_n755_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT110), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT111), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n578_), .A2(G85gat), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT112), .Z(new_n787_));
  AOI21_X1  g586(.A(new_n782_), .B1(new_n785_), .B2(new_n787_), .ZN(G1336gat));
  AOI21_X1  g587(.A(G92gat), .B1(new_n781_), .B2(new_n678_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n678_), .A2(G92gat), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT113), .Z(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n785_), .B2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT114), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n784_), .B2(new_n661_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n248_), .A2(new_n250_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n795_), .A3(new_n660_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  XOR2_X1   g597(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(G106gat), .B(new_n801_), .C1(new_n783_), .C2(new_n662_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n799_), .A2(new_n800_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n781_), .A2(new_n235_), .A3(new_n690_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n803_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT117), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(KEYINPUT117), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g610(.A(new_n365_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(KEYINPUT55), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n353_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n361_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(KEYINPUT55), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n374_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n818_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n376_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n402_), .B1(new_n384_), .B2(new_n395_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n393_), .A2(new_n394_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n404_), .A2(new_n409_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n305_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n376_), .A2(new_n377_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n823_), .A2(new_n413_), .B1(new_n835_), .B2(new_n827_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(new_n303_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n822_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n818_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n413_), .B(new_n372_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n827_), .A2(new_n835_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n291_), .A2(new_n295_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(KEYINPUT57), .A3(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n832_), .A2(new_n837_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n350_), .A2(new_n414_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n846_), .B2(new_n380_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n846_), .A2(new_n380_), .A3(KEYINPUT54), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n845_), .A2(new_n349_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n678_), .A2(new_n674_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n849_), .A2(new_n632_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n413_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n849_), .A2(new_n851_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n632_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n859_));
  NAND2_X1  g658(.A1(new_n852_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n414_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n853_), .B1(new_n861_), .B2(G113gat), .ZN(G1340gat));
  AOI21_X1  g661(.A(new_n379_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n845_), .A2(new_n349_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n848_), .A2(new_n847_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n522_), .B1(new_n379_), .B2(KEYINPUT60), .ZN(new_n867_));
  AND4_X1   g666(.A1(new_n855_), .A2(new_n866_), .A3(new_n850_), .A4(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n522_), .A2(KEYINPUT60), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n868_), .A2(KEYINPUT120), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT120), .B1(new_n868_), .B2(new_n870_), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n863_), .A2(new_n522_), .B1(new_n871_), .B2(new_n872_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n852_), .B2(new_n708_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n349_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G127gat), .ZN(G1342gat));
  XNOR2_X1  g675(.A(KEYINPUT122), .B(G134gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n305_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n879_));
  AOI211_X1 g678(.A(KEYINPUT121), .B(G134gat), .C1(new_n852_), .C2(new_n303_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n852_), .A2(new_n303_), .ZN(new_n882_));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n879_), .A2(new_n880_), .A3(new_n884_), .ZN(G1343gat));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  INV_X1    g685(.A(new_n626_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n854_), .B2(new_n887_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n849_), .A2(KEYINPUT123), .A3(new_n626_), .A4(new_n851_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n413_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G141gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n866_), .A2(new_n887_), .A3(new_n850_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT123), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n854_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n536_), .A3(new_n413_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n896_), .ZN(G1344gat));
  OAI21_X1  g696(.A(new_n380_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G148gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n537_), .A3(new_n380_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1345gat));
  OAI21_X1  g700(.A(new_n708_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT124), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n895_), .A2(new_n708_), .A3(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n895_), .B2(new_n303_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n305_), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n287_), .B(new_n910_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1347gat));
  NOR4_X1   g711(.A1(new_n849_), .A2(new_n578_), .A3(new_n632_), .A4(new_n680_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n399_), .B1(new_n913_), .B2(new_n413_), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT57), .B1(new_n842_), .B2(new_n843_), .ZN(new_n915_));
  AOI211_X1 g714(.A(new_n833_), .B(new_n303_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n708_), .B1(new_n917_), .B2(new_n832_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n865_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n674_), .B(new_n678_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n467_), .A2(new_n468_), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n920_), .A2(new_n414_), .A3(new_n632_), .A4(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n914_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(KEYINPUT62), .B2(new_n914_), .ZN(G1348gat));
  NAND2_X1  g723(.A1(new_n913_), .A2(new_n380_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n438_), .A2(new_n417_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n913_), .A2(new_n708_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT125), .ZN(new_n929_));
  INV_X1    g728(.A(new_n913_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n460_), .B1(new_n930_), .B2(new_n349_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n913_), .A2(new_n932_), .A3(new_n708_), .A4(new_n927_), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n929_), .A2(new_n931_), .A3(new_n933_), .ZN(G1350gat));
  OAI21_X1  g733(.A(G190gat), .B1(new_n930_), .B2(new_n910_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n303_), .B1(new_n440_), .B2(new_n439_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n930_), .B2(new_n936_), .ZN(G1351gat));
  NAND4_X1  g736(.A1(new_n866_), .A2(new_n674_), .A3(new_n887_), .A4(new_n678_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n414_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(G197gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n938_), .A2(new_n379_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n448_), .ZN(G1353gat));
  NOR4_X1   g742(.A1(new_n849_), .A2(new_n578_), .A3(new_n626_), .A4(new_n680_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945_));
  INV_X1    g744(.A(G211gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n944_), .A2(new_n708_), .A3(new_n947_), .A4(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n938_), .A2(new_n349_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n952_), .A2(KEYINPUT127), .A3(new_n947_), .A4(new_n948_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n945_), .B(new_n946_), .C1(new_n938_), .C2(new_n349_), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n951_), .A2(new_n953_), .A3(new_n954_), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n944_), .B2(new_n303_), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n305_), .A2(G218gat), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n944_), .B2(new_n957_), .ZN(G1355gat));
endmodule


