//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G8gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  INV_X1    g005(.A(G22gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G15gat), .A2(G22gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G1gat), .A2(G8gat), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n208_), .A2(new_n209_), .B1(KEYINPUT14), .B2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n205_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G29gat), .B(G36gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n217_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n222_), .A3(new_n213_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n202_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n220_), .A2(KEYINPUT15), .A3(new_n217_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n214_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT76), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n214_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n202_), .B(KEYINPUT77), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n224_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n235_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(new_n224_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n250_), .A3(KEYINPUT64), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n256_));
  INV_X1    g055(.A(G106gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(G85gat), .A3(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G85gat), .B(G92gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT9), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n255_), .A2(new_n259_), .A3(new_n261_), .A4(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n262_), .A2(KEYINPUT8), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT7), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT65), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n274_), .A3(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n267_), .B1(new_n255_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT8), .ZN(new_n278_));
  NOR4_X1   g077(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n251_), .B(new_n268_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n281_), .B2(new_n263_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n265_), .B(new_n222_), .C1(new_n277_), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G232gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT34), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n248_), .A2(new_n250_), .A3(KEYINPUT64), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT64), .B1(new_n248_), .B2(new_n250_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n259_), .B(new_n261_), .C1(new_n260_), .C2(new_n262_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n279_), .A2(new_n280_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n249_), .B1(G99gat), .B2(G106gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n268_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n263_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT8), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n268_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n266_), .B1(new_n291_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n293_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n226_), .A2(new_n227_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n283_), .B(new_n288_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n286_), .A2(new_n287_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n265_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n228_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n305_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n288_), .A4(new_n283_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT73), .A3(new_n310_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G190gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT36), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT37), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n306_), .A2(new_n310_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n311_), .A2(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n324_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n328_), .B2(KEYINPUT37), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n306_), .A2(new_n310_), .A3(new_n323_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n318_), .B1(new_n306_), .B2(new_n310_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n326_), .B(KEYINPUT37), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n325_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT74), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(new_n325_), .C1(new_n329_), .C2(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G57gat), .B(G64gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G71gat), .B(G78gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT11), .ZN(new_n341_));
  XOR2_X1   g140(.A(G71gat), .B(G78gat), .Z(new_n342_));
  INV_X1    g141(.A(G64gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G57gat), .ZN(new_n344_));
  INV_X1    g143(.A(G57gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G64gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n346_), .A3(KEYINPUT11), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n339_), .A2(KEYINPUT11), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n341_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n214_), .B(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(G231gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G155gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT16), .ZN(new_n357_));
  XOR2_X1   g156(.A(G183gat), .B(G211gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT17), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n355_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(KEYINPUT17), .B2(new_n360_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n354_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT67), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n350_), .A2(new_n361_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT66), .B(new_n341_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT12), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n302_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT12), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n302_), .B2(new_n350_), .ZN(new_n373_));
  AND2_X1   g172(.A1(G230gat), .A2(G233gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n302_), .B2(new_n350_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n369_), .A2(KEYINPUT12), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n307_), .A2(KEYINPUT67), .A3(new_n368_), .A4(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n371_), .A2(new_n373_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n302_), .A2(new_n350_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n307_), .A2(new_n351_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G120gat), .B(G148gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT5), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G176gat), .B(G204gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT68), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n378_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT69), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(KEYINPUT13), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n394_));
  NAND3_X1  g193(.A1(new_n389_), .A2(new_n390_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n338_), .A2(new_n366_), .A3(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G211gat), .B(G218gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT84), .B(G204gat), .ZN(new_n399_));
  INV_X1    g198(.A(G197gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT21), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(G197gat), .B2(G204gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n398_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n407_), .B2(KEYINPUT21), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT85), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(KEYINPUT21), .A3(new_n398_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT25), .B(G183gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT26), .B(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G169gat), .ZN(new_n415_));
  INV_X1    g214(.A(G176gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT24), .A3(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n417_), .A2(KEYINPUT24), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G183gat), .ZN(new_n423_));
  INV_X1    g222(.A(G190gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT23), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT23), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(G183gat), .A3(G190gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n426_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n418_), .A2(KEYINPUT88), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n418_), .A2(KEYINPUT88), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G169gat), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n432_), .B(new_n433_), .C1(new_n416_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n425_), .A2(new_n427_), .A3(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT78), .B(KEYINPUT23), .C1(new_n423_), .C2(new_n424_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n437_), .B(new_n438_), .C1(G183gat), .C2(G190gat), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n422_), .A2(new_n431_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n411_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT19), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT20), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n409_), .A2(new_n410_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n431_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(new_n415_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n437_), .A2(new_n438_), .ZN(new_n451_));
  OAI22_X1  g250(.A1(new_n448_), .A2(new_n450_), .B1(new_n421_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n445_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n441_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT89), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n411_), .A2(new_n440_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT20), .B1(new_n446_), .B2(new_n452_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n443_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT18), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G64gat), .B(G92gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n454_), .A2(KEYINPUT89), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n441_), .B2(new_n453_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n458_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n462_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT96), .B(KEYINPUT27), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT27), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n446_), .A2(new_n452_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n441_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n443_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n456_), .A2(new_n457_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(new_n443_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n473_), .B1(new_n479_), .B2(new_n468_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n463_), .A3(KEYINPUT95), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT95), .B1(new_n480_), .B2(new_n463_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n472_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT3), .Z(new_n490_));
  NAND2_X1  g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n491_), .B(KEYINPUT2), .Z(new_n492_));
  OAI211_X1 g291(.A(new_n487_), .B(new_n488_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT1), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n488_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n487_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n489_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n491_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n411_), .B1(KEYINPUT29), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(KEYINPUT86), .A2(G228gat), .A3(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT86), .B1(G228gat), .B2(G233gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT87), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n499_), .A2(KEYINPUT29), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT28), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G22gat), .B(G50gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n510_), .A2(KEYINPUT28), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(KEYINPUT28), .ZN(new_n515_));
  INV_X1    g314(.A(new_n512_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n509_), .B1(new_n513_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n508_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n520_), .A3(new_n517_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n507_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n513_), .A2(new_n520_), .A3(new_n517_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n505_), .B(new_n506_), .C1(new_n523_), .C2(new_n518_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT82), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G120gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(new_n499_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n499_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G225gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(KEYINPUT90), .A3(KEYINPUT4), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n532_), .A2(KEYINPUT4), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n531_), .A2(KEYINPUT4), .A3(new_n532_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n542_), .B2(new_n535_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G29gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G85gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT0), .B(G57gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n534_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n550_), .B2(new_n536_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G227gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT81), .ZN(new_n555_));
  XOR2_X1   g354(.A(G71gat), .B(G99gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n452_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n530_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G15gat), .B(G43gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT80), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT30), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT31), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n559_), .B(new_n563_), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n553_), .A2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n484_), .A2(new_n526_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n467_), .B2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n455_), .A2(KEYINPUT93), .A3(new_n458_), .A4(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n479_), .A2(new_n569_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n552_), .A2(new_n570_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(KEYINPUT91), .A2(KEYINPUT33), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n551_), .A2(new_n574_), .ZN(new_n575_));
  OAI221_X1 g374(.A(new_n547_), .B1(KEYINPUT91), .B2(KEYINPUT33), .C1(new_n550_), .C2(new_n536_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n547_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n542_), .B2(new_n535_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT92), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n577_), .C1(new_n542_), .C2(new_n535_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n575_), .A2(new_n576_), .A3(new_n579_), .A4(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n573_), .B1(new_n470_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n525_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n525_), .A2(new_n552_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n585_), .B(new_n472_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n564_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n566_), .B1(new_n587_), .B2(KEYINPUT97), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589_));
  INV_X1    g388(.A(new_n483_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n590_), .A2(new_n481_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n591_), .A2(new_n585_), .B1(new_n583_), .B2(new_n525_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n592_), .B2(new_n564_), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n246_), .B(new_n397_), .C1(new_n588_), .C2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G1gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n552_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT99), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n320_), .A2(new_n324_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n396_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n366_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n603_), .A2(new_n246_), .A3(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(new_n552_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n596_), .A2(new_n597_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT98), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(KEYINPUT98), .ZN(new_n610_));
  OAI221_X1 g409(.A(new_n599_), .B1(new_n595_), .B2(new_n607_), .C1(new_n609_), .C2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(G8gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n594_), .A2(new_n612_), .A3(new_n484_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n602_), .A2(new_n484_), .A3(new_n605_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n616_));
  AND4_X1   g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .A4(G8gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n612_), .B1(KEYINPUT100), .B2(KEYINPUT39), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n615_), .A2(new_n618_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT102), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n622_), .B(new_n613_), .C1(new_n617_), .C2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n621_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  AOI21_X1  g428(.A(new_n206_), .B1(new_n606_), .B2(new_n564_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n594_), .A2(new_n206_), .A3(new_n564_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  AOI21_X1  g432(.A(new_n207_), .B1(new_n606_), .B2(new_n526_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT42), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n594_), .A2(new_n207_), .A3(new_n526_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1327gat));
  NOR3_X1   g436(.A1(new_n603_), .A2(new_n246_), .A3(new_n366_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n588_), .A2(new_n593_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n337_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT37), .B1(new_n330_), .B2(new_n331_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT72), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n332_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n336_), .B1(new_n644_), .B2(new_n325_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n639_), .B1(new_n640_), .B2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT43), .B(new_n338_), .C1(new_n588_), .C2(new_n593_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n638_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT44), .B(new_n638_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n552_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n246_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n604_), .A2(new_n601_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n603_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n553_), .A2(G29gat), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT103), .Z(new_n661_));
  OAI21_X1  g460(.A(new_n655_), .B1(new_n659_), .B2(new_n661_), .ZN(G1328gat));
  NAND2_X1  g461(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n663_));
  NOR2_X1   g462(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT105), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n651_), .A2(new_n484_), .A3(new_n652_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n591_), .A2(G36gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n659_), .B2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n656_), .A2(KEYINPUT45), .A3(new_n658_), .A4(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n663_), .B(new_n665_), .C1(new_n667_), .C2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n665_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n666_), .B2(G36gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n663_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n674_), .A2(new_n678_), .ZN(G1329gat));
  NAND4_X1  g478(.A1(new_n651_), .A2(G43gat), .A3(new_n564_), .A4(new_n652_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n564_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n659_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(G43gat), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1330gat));
  OR3_X1    g484(.A1(new_n659_), .A2(G50gat), .A3(new_n525_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n653_), .A2(KEYINPUT107), .A3(new_n526_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G50gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT107), .B1(new_n653_), .B2(new_n526_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n603_), .A2(new_n246_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n604_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n602_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n553_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n245_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n646_), .A2(new_n604_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n603_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n345_), .A3(new_n552_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n699_), .ZN(G1332gat));
  AOI21_X1  g499(.A(new_n343_), .B1(new_n693_), .B2(new_n484_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT48), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n343_), .A3(new_n484_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1333gat));
  INV_X1    g503(.A(G71gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n693_), .B2(new_n564_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT49), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(new_n705_), .A3(new_n564_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1334gat));
  INV_X1    g508(.A(G78gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n693_), .B2(new_n526_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT50), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n698_), .A2(new_n710_), .A3(new_n526_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1335gat));
  OR2_X1    g513(.A1(new_n647_), .A2(new_n648_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n691_), .A2(new_n366_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n553_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n657_), .A2(new_n396_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n696_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n553_), .A2(G85gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1336gat));
  NAND2_X1  g522(.A1(new_n484_), .A2(G92gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT108), .Z(new_n725_));
  NOR2_X1   g524(.A1(new_n721_), .A2(new_n591_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n717_), .A2(new_n725_), .B1(new_n726_), .B2(G92gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT109), .ZN(G1337gat));
  OAI21_X1  g527(.A(G99gat), .B1(new_n717_), .B2(new_n681_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n720_), .A2(new_n564_), .A3(new_n256_), .A4(new_n258_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g531(.A(new_n526_), .B(new_n716_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G106gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n733_), .A2(KEYINPUT110), .A3(G106gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(KEYINPUT52), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT110), .B1(new_n733_), .B2(G106gat), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n525_), .A2(G106gat), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n739_), .A2(new_n740_), .B1(new_n720_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT53), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n738_), .A2(new_n742_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1339gat));
  NOR4_X1   g546(.A1(new_n484_), .A2(new_n681_), .A3(new_n526_), .A4(new_n553_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  INV_X1    g549(.A(new_n223_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n234_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n233_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n221_), .A2(new_n223_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n240_), .B1(new_n754_), .B2(new_n234_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n241_), .A2(new_n390_), .A3(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n302_), .A2(new_n370_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n758_), .A2(KEYINPUT67), .B1(new_n380_), .B2(new_n372_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n759_), .A2(KEYINPUT55), .A3(new_n371_), .A4(new_n375_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n378_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n371_), .A2(new_n373_), .A3(new_n379_), .A4(new_n377_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n374_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n388_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n388_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n757_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n750_), .B1(new_n646_), .B2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(new_n335_), .A3(new_n750_), .A4(new_n337_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n768_), .A2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n245_), .B(new_n390_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n391_), .A2(new_n241_), .A3(new_n756_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n600_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(KEYINPUT111), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n601_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT57), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n604_), .B1(new_n775_), .B2(new_n786_), .ZN(new_n787_));
  OR3_X1    g586(.A1(new_n397_), .A2(KEYINPUT54), .A3(new_n245_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT54), .B1(new_n397_), .B2(new_n245_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n749_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G113gat), .B1(new_n791_), .B2(new_n245_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n790_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n779_), .A2(new_n780_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT114), .B(new_n794_), .C1(new_n771_), .C2(new_n774_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n785_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n793_), .B1(new_n799_), .B2(new_n604_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n749_), .A2(KEYINPUT59), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n795_), .A2(new_n796_), .B1(KEYINPUT57), .B2(new_n783_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n366_), .B1(new_n805_), .B2(new_n798_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n804_), .B(new_n801_), .C1(new_n806_), .C2(new_n793_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n787_), .A2(new_n790_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n748_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(KEYINPUT59), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n809_), .A2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n246_), .A2(KEYINPUT116), .ZN(new_n819_));
  MUX2_X1   g618(.A(KEYINPUT116), .B(new_n819_), .S(G113gat), .Z(new_n820_));
  AOI21_X1  g619(.A(new_n792_), .B1(new_n818_), .B2(new_n820_), .ZN(G1340gat));
  AOI21_X1  g620(.A(new_n396_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n808_), .A2(KEYINPUT117), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT117), .B1(new_n808_), .B2(new_n822_), .ZN(new_n824_));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n396_), .B2(KEYINPUT60), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n825_), .A2(KEYINPUT60), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n791_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT118), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n808_), .A2(new_n822_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G120gat), .B1(new_n833_), .B2(KEYINPUT117), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n832_), .B(new_n829_), .C1(new_n834_), .C2(new_n823_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(G1341gat));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n791_), .A2(new_n837_), .A3(new_n366_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n809_), .A2(new_n604_), .A3(new_n817_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g639(.A(G134gat), .B1(new_n791_), .B2(new_n601_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT119), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n646_), .A2(G134gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n818_), .B2(new_n843_), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n564_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n591_), .A2(new_n526_), .A3(new_n552_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n245_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n848_), .A2(new_n396_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT120), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NAND2_X1  g653(.A1(new_n849_), .A2(new_n366_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT121), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT61), .B(G155gat), .Z(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  AOI21_X1  g657(.A(G162gat), .B1(new_n849_), .B2(new_n601_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n646_), .A2(G162gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT122), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n849_), .B2(new_n861_), .ZN(G1347gat));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  INV_X1    g662(.A(new_n800_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n591_), .A2(new_n565_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n525_), .B1(new_n865_), .B2(KEYINPUT123), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(KEYINPUT123), .B2(new_n865_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n246_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n863_), .B1(new_n869_), .B2(new_n415_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n434_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT62), .B(G169gat), .C1(new_n868_), .C2(new_n246_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1348gat));
  AND2_X1   g674(.A1(new_n867_), .A2(new_n810_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(G176gat), .A3(new_n603_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT125), .Z(new_n878_));
  INV_X1    g677(.A(new_n868_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G176gat), .B1(new_n879_), .B2(new_n603_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1349gat));
  AOI21_X1  g680(.A(G183gat), .B1(new_n876_), .B2(new_n366_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n604_), .A2(new_n412_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n879_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n868_), .B2(new_n338_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n601_), .A2(new_n413_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n868_), .B2(new_n886_), .ZN(G1351gat));
  AND2_X1   g686(.A1(new_n484_), .A2(new_n585_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n845_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n246_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n400_), .ZN(G1352gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n396_), .ZN(new_n892_));
  MUX2_X1   g691(.A(G204gat), .B(new_n399_), .S(new_n892_), .Z(G1353gat));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n604_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n894_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(G1354gat));
  INV_X1    g699(.A(new_n889_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G218gat), .B1(new_n901_), .B2(new_n601_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n646_), .A2(G218gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT127), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n901_), .B2(new_n904_), .ZN(G1355gat));
endmodule


