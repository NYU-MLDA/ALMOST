//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204_));
  AND2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT1), .ZN(new_n207_));
  OR2_X1    g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n204_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n210_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n216_), .A2(new_n219_), .A3(KEYINPUT88), .A4(new_n209_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(KEYINPUT2), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n210_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n225_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n205_), .A2(new_n206_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n221_), .A2(new_n222_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n222_), .B1(new_n221_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n203_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n234_), .B(KEYINPUT93), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G78gat), .B(G106gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n239_));
  AND2_X1   g038(.A1(G197gat), .A2(G204gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT21), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  INV_X1    g044(.A(G218gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n246_), .A2(G211gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(G211gat), .ZN(new_n248_));
  OAI22_X1  g047(.A1(new_n247_), .A2(new_n248_), .B1(new_n241_), .B2(new_n240_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n244_), .B1(new_n250_), .B2(KEYINPUT21), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n212_), .A2(new_n220_), .B1(new_n230_), .B2(new_n229_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n203_), .ZN(new_n253_));
  INV_X1    g052(.A(G233gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G228gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(G228gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n221_), .A2(new_n231_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT89), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n252_), .A2(new_n222_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(KEYINPUT29), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n251_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI221_X4 g065(.A(new_n238_), .B1(new_n253_), .B2(new_n259_), .C1(new_n263_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n266_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n253_), .A2(new_n259_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n237_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT28), .B(G22gat), .ZN(new_n271_));
  INV_X1    g070(.A(G50gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT90), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n267_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n232_), .A2(new_n233_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n265_), .B1(new_n277_), .B2(KEYINPUT29), .ZN(new_n278_));
  INV_X1    g077(.A(new_n269_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n238_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n268_), .A2(new_n269_), .A3(new_n237_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n276_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n236_), .B1(new_n275_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n274_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n281_), .A3(new_n276_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n235_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G127gat), .B(G134gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n261_), .A2(new_n289_), .A3(new_n262_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n260_), .A2(new_n289_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT4), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n261_), .A2(new_n293_), .A3(new_n289_), .A4(new_n262_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT97), .Z(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n290_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G85gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G57gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n283_), .A2(new_n286_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT19), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n251_), .ZN(new_n312_));
  INV_X1    g111(.A(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n315_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n323_));
  AND2_X1   g122(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n323_), .B(KEYINPUT22), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327_));
  AOI21_X1  g126(.A(G176gat), .B1(new_n327_), .B2(G169gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT83), .B(G169gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n323_), .B1(new_n330_), .B2(KEYINPUT22), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n322_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT25), .B(G183gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT26), .B(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(G169gat), .B2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n313_), .A2(new_n314_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n333_), .A2(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT82), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n339_), .A2(new_n342_), .A3(new_n346_), .A4(new_n343_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n338_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n332_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n332_), .A2(new_n348_), .A3(KEYINPUT85), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n312_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n344_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n338_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n314_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n342_), .A2(new_n321_), .A3(new_n343_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n357_), .B(new_n358_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n355_), .B(new_n359_), .C1(new_n361_), .C2(new_n244_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT20), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n311_), .B1(new_n353_), .B2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n351_), .A2(new_n352_), .A3(new_n312_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n355_), .A2(new_n359_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n251_), .A2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n367_), .A2(KEYINPUT20), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n368_), .A3(new_n310_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G8gat), .B(G36gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT100), .B1(new_n370_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT100), .ZN(new_n377_));
  INV_X1    g176(.A(new_n375_), .ZN(new_n378_));
  AOI211_X1 g177(.A(new_n377_), .B(new_n378_), .C1(new_n364_), .C2(new_n369_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT27), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n332_), .A2(new_n348_), .A3(KEYINPUT85), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT85), .B1(new_n332_), .B2(new_n348_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n251_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT94), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n355_), .A2(new_n359_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n312_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n310_), .A2(KEYINPUT20), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n362_), .B2(KEYINPUT94), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n367_), .A2(KEYINPUT20), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n381_), .A2(new_n382_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n312_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n389_), .B(new_n378_), .C1(new_n392_), .C2(new_n310_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT101), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n380_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n308_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n386_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(new_n353_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n310_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n375_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(KEYINPUT96), .A3(new_n393_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n389_), .B1(new_n392_), .B2(new_n310_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n375_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT102), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n401_), .A2(KEYINPUT102), .A3(new_n402_), .A4(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n283_), .A2(new_n286_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n378_), .A2(KEYINPUT32), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n403_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n370_), .A2(new_n412_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n413_), .B(new_n414_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n401_), .A2(new_n405_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n290_), .A2(KEYINPUT4), .A3(new_n291_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n294_), .A2(new_n295_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT99), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT99), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n292_), .A2(new_n420_), .A3(new_n295_), .A4(new_n294_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n290_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT98), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n302_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n422_), .B2(new_n302_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n419_), .B(new_n421_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n304_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n297_), .A2(KEYINPUT33), .A3(new_n298_), .A4(new_n303_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n415_), .B1(new_n416_), .B2(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n396_), .A2(new_n410_), .B1(new_n411_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G43gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n434_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n391_), .B(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT87), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(KEYINPUT87), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n438_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n438_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n289_), .B(KEYINPUT31), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n202_), .B1(new_n432_), .B2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n284_), .A2(new_n235_), .A3(new_n285_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n235_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n297_), .A2(new_n298_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n302_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n304_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n380_), .A2(new_n394_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n410_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n431_), .A2(new_n411_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n450_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(KEYINPUT103), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n456_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n395_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n411_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n451_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT67), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(G99gat), .ZN(new_n473_));
  INV_X1    g272(.A(G106gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT6), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n469_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n472_), .A2(new_n478_), .A3(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G85gat), .B(G92gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(KEYINPUT68), .A3(new_n484_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT8), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n480_), .A2(new_n469_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n478_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n475_), .A2(KEYINPUT64), .A3(new_n477_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT65), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(KEYINPUT65), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n484_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT66), .B1(new_n494_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n490_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n493_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT64), .B1(new_n475_), .B2(new_n477_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n499_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n500_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n502_), .A2(new_n503_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT10), .B(G99gat), .Z(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n474_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n484_), .A2(KEYINPUT9), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT9), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n489_), .A2(new_n508_), .B1(new_n510_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n522_));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n519_), .A2(new_n526_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n468_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n489_), .A2(new_n508_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT69), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n510_), .A2(new_n518_), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT69), .B1(new_n509_), .B2(new_n517_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n524_), .A2(KEYINPUT12), .A3(new_n525_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n527_), .C1(new_n529_), .C2(KEYINPUT12), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n530_), .B1(new_n540_), .B2(new_n468_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G120gat), .B(G148gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT71), .ZN(new_n543_));
  XOR2_X1   g342(.A(G176gat), .B(G204gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n541_), .B(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n541_), .A2(new_n548_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n541_), .A2(new_n548_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n556_), .B(new_n557_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G29gat), .B(G36gat), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT73), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT73), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT15), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572_));
  INV_X1    g371(.A(G1gat), .ZN(new_n573_));
  INV_X1    g372(.A(G8gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G1gat), .B(G8gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT79), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n581_), .B(new_n582_), .C1(new_n578_), .C2(new_n569_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n569_), .B(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(G229gat), .A3(G233gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT81), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT80), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n586_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n592_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n560_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n467_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n533_), .A2(new_n534_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n508_), .B2(new_n489_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n569_), .B(KEYINPUT15), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT74), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n536_), .A2(new_n603_), .A3(new_n571_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n510_), .A2(new_n518_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n569_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n531_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT75), .B1(new_n519_), .B2(new_n606_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n602_), .B(new_n604_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT34), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT35), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(KEYINPUT36), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n613_), .B(KEYINPUT35), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n536_), .B2(new_n571_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n621_), .B(KEYINPUT76), .C1(new_n609_), .C2(new_n610_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n607_), .A2(new_n608_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n519_), .A2(KEYINPUT75), .A3(new_n606_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT76), .B1(new_n626_), .B2(new_n621_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n615_), .B(new_n619_), .C1(new_n623_), .C2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n618_), .B(KEYINPUT36), .Z(new_n629_));
  OAI21_X1  g428(.A(new_n621_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT76), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n632_), .A2(new_n622_), .B1(new_n614_), .B2(new_n611_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT77), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n615_), .B(new_n634_), .C1(new_n623_), .C2(new_n627_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n598_), .B(new_n628_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT78), .ZN(new_n639_));
  INV_X1    g438(.A(new_n629_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n628_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n641_), .B2(KEYINPUT37), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n615_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT77), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n636_), .A3(new_n629_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n639_), .A3(new_n598_), .A4(new_n628_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n526_), .B(new_n578_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT17), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G127gat), .B(G155gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT16), .ZN(new_n654_));
  XOR2_X1   g453(.A(G183gat), .B(G211gat), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n651_), .A2(new_n652_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(KEYINPUT17), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n648_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n597_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n573_), .A3(new_n456_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n450_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n466_), .B1(new_n666_), .B2(KEYINPUT103), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n432_), .A2(new_n202_), .A3(new_n450_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n646_), .A2(new_n628_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n560_), .A2(new_n660_), .A3(new_n595_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n307_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n663_), .A2(new_n664_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n665_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT104), .ZN(G1324gat));
  INV_X1    g477(.A(new_n465_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n662_), .A2(new_n574_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  INV_X1    g480(.A(new_n674_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n679_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(G8gat), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT39), .B(new_n574_), .C1(new_n682_), .C2(new_n679_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n674_), .B2(new_n462_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n662_), .A2(new_n436_), .A3(new_n450_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT106), .Z(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n674_), .B2(new_n411_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  INV_X1    g496(.A(G22gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n411_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n662_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1327gat));
  NOR2_X1   g500(.A1(new_n670_), .A2(new_n659_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n597_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n456_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n648_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT43), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n708_), .B(new_n648_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n593_), .A2(new_n594_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n559_), .A2(new_n660_), .A3(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT107), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(KEYINPUT108), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n709_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n708_), .B1(new_n467_), .B2(new_n648_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n713_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n710_), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n713_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n714_), .A2(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n456_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n705_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  INV_X1    g526(.A(G36gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n724_), .B2(new_n679_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n465_), .B(KEYINPUT110), .Z(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n704_), .A2(new_n728_), .A3(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT45), .Z(new_n733_));
  OAI21_X1  g532(.A(new_n727_), .B1(new_n729_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n719_), .A2(new_n714_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n722_), .A2(new_n723_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n679_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G36gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n732_), .B(KEYINPUT45), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(KEYINPUT46), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n734_), .A2(new_n740_), .ZN(G1329gat));
  NAND4_X1  g540(.A1(new_n735_), .A2(new_n736_), .A3(G43gat), .A4(new_n450_), .ZN(new_n742_));
  INV_X1    g541(.A(G43gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n703_), .B2(new_n462_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT47), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n272_), .B1(new_n724_), .B2(new_n699_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n699_), .A2(new_n272_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT111), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n704_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n735_), .A2(new_n699_), .A3(new_n736_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G50gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT112), .A3(new_n754_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1331gat));
  NOR2_X1   g559(.A1(new_n669_), .A2(new_n711_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n761_), .A2(new_n661_), .A3(new_n560_), .ZN(new_n762_));
  INV_X1    g561(.A(G57gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n456_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n672_), .A2(new_n659_), .A3(new_n595_), .A4(new_n560_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n307_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT113), .Z(G1332gat));
  OAI21_X1  g567(.A(G64gat), .B1(new_n765_), .B2(new_n730_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT48), .ZN(new_n770_));
  INV_X1    g569(.A(G64gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n771_), .A3(new_n731_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n765_), .B2(new_n462_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n762_), .A2(new_n776_), .A3(new_n450_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1334gat));
  OAI21_X1  g577(.A(G78gat), .B1(new_n765_), .B2(new_n411_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT50), .ZN(new_n780_));
  INV_X1    g579(.A(G78gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n762_), .A2(new_n781_), .A3(new_n699_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n711_), .A2(new_n659_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n710_), .A2(new_n560_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n307_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n761_), .A2(new_n560_), .A3(new_n702_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n514_), .A3(new_n456_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(G1336gat));
  OAI21_X1  g591(.A(G92gat), .B1(new_n786_), .B2(new_n730_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n515_), .A3(new_n679_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n790_), .A2(new_n511_), .A3(new_n450_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n786_), .A2(new_n462_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n473_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT51), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n796_), .B(new_n800_), .C1(new_n797_), .C2(new_n473_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n790_), .A2(new_n474_), .A3(new_n699_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n710_), .A2(new_n699_), .A3(new_n560_), .A4(new_n784_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(G106gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(G106gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT53), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n803_), .B(new_n810_), .C1(new_n807_), .C2(new_n806_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n540_), .B2(new_n468_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n540_), .A2(new_n468_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n815_), .A2(new_n816_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n540_), .A2(new_n814_), .A3(new_n468_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n548_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n555_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n578_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n582_), .B1(new_n606_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n581_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n590_), .B1(new_n584_), .B2(new_n582_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n586_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n590_), .B2(new_n833_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n824_), .A2(new_n711_), .B1(new_n549_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n813_), .B1(new_n835_), .B2(new_n671_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n548_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n821_), .A2(new_n822_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n711_), .B(new_n556_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n549_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT57), .A3(new_n670_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n583_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n843_));
  OR2_X1    g642(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n843_), .B(new_n844_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n556_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n824_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n834_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n648_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n836_), .A2(new_n842_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n660_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT54), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n595_), .A2(new_n659_), .A3(new_n855_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(new_n560_), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n857_), .A2(new_n648_), .B1(new_n854_), .B2(KEYINPUT54), .ZN(new_n858_));
  INV_X1    g657(.A(new_n648_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n560_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n854_), .A2(KEYINPUT54), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n853_), .A2(new_n863_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n679_), .A2(new_n462_), .A3(new_n699_), .A4(new_n307_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n595_), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n867_), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT118), .B1(new_n867_), .B2(G113gat), .ZN(new_n869_));
  INV_X1    g668(.A(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT59), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n866_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n711_), .A2(G113gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT119), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n868_), .A2(new_n869_), .B1(new_n874_), .B2(new_n876_), .ZN(G1340gat));
  AOI21_X1  g676(.A(new_n559_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n559_), .A2(KEYINPUT60), .ZN(new_n881_));
  MUX2_X1   g680(.A(KEYINPUT60), .B(new_n881_), .S(new_n879_), .Z(new_n882_));
  AND3_X1   g681(.A1(new_n870_), .A2(new_n880_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n880_), .B1(new_n870_), .B2(new_n882_), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n878_), .A2(new_n879_), .B1(new_n883_), .B2(new_n884_), .ZN(G1341gat));
  AOI21_X1  g684(.A(G127gat), .B1(new_n870_), .B2(new_n659_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(G127gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n659_), .A2(KEYINPUT121), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(G127gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n874_), .B2(new_n890_), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n870_), .A2(new_n892_), .A3(new_n671_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n859_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n892_), .ZN(G1343gat));
  AOI21_X1  g694(.A(new_n450_), .B1(new_n853_), .B2(new_n863_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n731_), .A2(new_n411_), .A3(new_n307_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(KEYINPUT122), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n896_), .B2(new_n897_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n711_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT123), .B(G141gat), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n711_), .B(new_n902_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1344gat));
  OAI21_X1  g705(.A(new_n560_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G148gat), .ZN(new_n908_));
  INV_X1    g707(.A(G148gat), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n909_), .B(new_n560_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1345gat));
  OAI21_X1  g710(.A(new_n659_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT61), .B(G155gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n913_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n659_), .B(new_n915_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1346gat));
  INV_X1    g716(.A(G162gat), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n918_), .B(new_n671_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n900_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n859_), .B1(new_n920_), .B2(new_n898_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n921_), .B2(new_n918_), .ZN(G1347gat));
  NAND3_X1  g721(.A1(new_n731_), .A2(new_n411_), .A3(new_n464_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n853_), .B2(new_n863_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n711_), .A2(new_n356_), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT124), .Z(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n313_), .B1(new_n924_), .B2(new_n711_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n929_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n927_), .B1(new_n930_), .B2(new_n931_), .ZN(G1348gat));
  NAND2_X1  g731(.A1(new_n924_), .A2(new_n560_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g733(.A1(new_n924_), .A2(new_n659_), .ZN(new_n935_));
  OR3_X1    g734(.A1(new_n935_), .A2(KEYINPUT125), .A3(new_n333_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(new_n935_), .B2(new_n333_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n319_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n924_), .A2(new_n671_), .A3(new_n334_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n924_), .A2(new_n648_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n320_), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n730_), .A2(new_n308_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n896_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n711_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n864_), .A2(new_n462_), .A3(new_n560_), .A4(new_n943_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(G204gat), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n896_), .A2(new_n950_), .A3(new_n560_), .A4(new_n943_), .ZN(new_n951_));
  INV_X1    g750(.A(G204gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n948_), .B2(KEYINPUT126), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n949_), .B1(new_n951_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n948_), .A2(KEYINPUT126), .ZN(new_n955_));
  AND4_X1   g754(.A1(KEYINPUT127), .A2(new_n955_), .A3(G204gat), .A4(new_n951_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n954_), .A2(new_n956_), .ZN(G1353gat));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  AND2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n944_), .B(new_n659_), .C1(new_n958_), .C2(new_n959_), .ZN(new_n960_));
  AND2_X1   g759(.A1(new_n944_), .A2(new_n659_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n958_), .ZN(G1354gat));
  NAND3_X1  g761(.A1(new_n944_), .A2(new_n246_), .A3(new_n671_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n944_), .A2(new_n648_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n246_), .ZN(G1355gat));
endmodule


