//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(new_n218_), .C1(G99gat), .C2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n210_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT66), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT66), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n213_), .B(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(KEYINPUT8), .C1(new_n226_), .C2(new_n206_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n204_), .A2(new_n228_), .A3(new_n205_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n219_), .A2(new_n221_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n214_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AOI211_X1 g032(.A(KEYINPUT65), .B(new_n229_), .C1(new_n214_), .C2(new_n230_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n223_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT66), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n214_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n207_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n216_), .B1(new_n240_), .B2(KEYINPUT8), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n215_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G29gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G232gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT34), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT35), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT8), .B1(new_n226_), .B2(new_n206_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT67), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n227_), .A3(new_n235_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n215_), .A3(new_n245_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n248_), .A2(new_n253_), .A3(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n251_), .A2(new_n252_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n259_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n261_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT74), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n260_), .A2(KEYINPUT74), .A3(new_n261_), .A4(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n260_), .A2(new_n261_), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n264_), .B(KEYINPUT36), .Z(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(KEYINPUT75), .A3(new_n273_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n271_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT37), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n278_), .A2(new_n279_), .B1(new_n271_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT79), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G15gat), .B(G22gat), .ZN(new_n283_));
  INV_X1    g082(.A(G1gat), .ZN(new_n284_));
  INV_X1    g083(.A(G8gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n283_), .B1(new_n286_), .B2(KEYINPUT76), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(KEYINPUT76), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G8gat), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT77), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G231gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT68), .B(G71gat), .ZN(new_n296_));
  INV_X1    g095(.A(G78gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n299_), .B(KEYINPUT11), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n295_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G155gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT17), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n295_), .A2(new_n304_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n311_), .A2(KEYINPUT17), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n305_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n305_), .A2(new_n313_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n282_), .B(new_n315_), .C1(new_n316_), .C2(new_n312_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n315_), .A2(new_n282_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n281_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT80), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT25), .B(G183gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT24), .A3(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n325_), .A2(KEYINPUT24), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT23), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(G183gat), .A3(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n337_));
  AOI21_X1  g136(.A(G176gat), .B1(new_n337_), .B2(KEYINPUT22), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n332_), .A2(new_n334_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(new_n340_), .B2(new_n334_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n339_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT86), .B(G43gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G15gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G71gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n349_), .B(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT87), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT31), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G99gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n353_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n349_), .B(new_n352_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n362_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G22gat), .B(G50gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G197gat), .ZN(new_n370_));
  INV_X1    g169(.A(G204gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(KEYINPUT21), .A3(new_n373_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n376_), .A2(KEYINPUT92), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n379_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT93), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n396_), .B(new_n397_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n389_), .B(new_n390_), .C1(new_n393_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(G155gat), .A3(G162gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT89), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n389_), .A2(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n404_), .A2(new_n405_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n399_), .B1(new_n394_), .B2(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(KEYINPUT88), .A2(G141gat), .A3(G148gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n401_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n385_), .B(new_n387_), .C1(new_n388_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n387_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n388_), .B1(new_n401_), .B2(new_n413_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n384_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n369_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n401_), .A2(new_n413_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n421_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT28), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT91), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n424_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(new_n422_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n415_), .A2(new_n418_), .A3(new_n369_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n420_), .A2(new_n428_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n428_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n419_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT19), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n384_), .A2(new_n336_), .A3(new_n344_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n342_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT22), .B(G169gat), .ZN(new_n442_));
  INV_X1    g241(.A(G176gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n326_), .A2(KEYINPUT94), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n326_), .A2(KEYINPUT94), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n335_), .B1(G183gat), .B2(G190gat), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n330_), .A2(new_n441_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT20), .B1(new_n449_), .B2(new_n384_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n439_), .B1(new_n440_), .B2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G8gat), .B(G36gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n385_), .A2(new_n345_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n449_), .B2(new_n384_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n439_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n455_), .B1(new_n451_), .B2(new_n460_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n437_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n440_), .A2(new_n450_), .A3(new_n439_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT99), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n456_), .A2(new_n458_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n439_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT99), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n455_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n461_), .A2(KEYINPUT27), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n464_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G29gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G85gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT0), .B(G57gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n401_), .A2(new_n413_), .A3(new_n356_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n357_), .A2(new_n359_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n414_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT95), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n421_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n484_), .A4(new_n481_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n483_), .A2(KEYINPUT4), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n484_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n480_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n487_), .B2(new_n481_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT4), .B1(new_n360_), .B2(new_n421_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n485_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n498_), .A2(new_n479_), .A3(new_n486_), .A4(new_n489_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n367_), .A2(new_n436_), .A3(new_n475_), .A4(new_n501_), .ZN(new_n502_));
  AND4_X1   g301(.A1(new_n432_), .A2(new_n495_), .A3(new_n435_), .A4(new_n499_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n473_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n440_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n450_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n459_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n470_), .B1(new_n507_), .B2(new_n469_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n466_), .A2(KEYINPUT99), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n510_), .B2(new_n455_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT100), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n503_), .A2(new_n511_), .A3(new_n512_), .A4(new_n464_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n495_), .A2(new_n432_), .A3(new_n435_), .A4(new_n499_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT100), .B1(new_n474_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n483_), .A2(KEYINPUT97), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT97), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n487_), .A2(new_n518_), .A3(new_n481_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n485_), .A3(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n484_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n480_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n522_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n499_), .A2(new_n524_), .A3(KEYINPUT33), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT33), .B1(new_n499_), .B2(new_n524_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT98), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT98), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n523_), .B(new_n529_), .C1(new_n526_), .C2(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n455_), .A2(KEYINPUT32), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n451_), .A2(new_n460_), .A3(new_n531_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n500_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n528_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n516_), .B1(new_n537_), .B2(new_n436_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n502_), .B1(new_n538_), .B2(new_n367_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G120gat), .B(G148gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT5), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G176gat), .B(G204gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT70), .ZN(new_n545_));
  INV_X1    g344(.A(G230gat), .ZN(new_n546_));
  INV_X1    g345(.A(G233gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n242_), .A2(new_n304_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n303_), .B(new_n215_), .C1(new_n236_), .C2(new_n241_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT12), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n242_), .A2(new_n552_), .A3(new_n304_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n548_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n548_), .B1(new_n550_), .B2(KEYINPUT69), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT69), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n242_), .B2(new_n304_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n550_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n545_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n548_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n550_), .A2(KEYINPUT12), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n303_), .B1(new_n256_), .B2(new_n215_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n553_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n560_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n555_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n557_), .A2(new_n550_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n544_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n559_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n559_), .B2(new_n570_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n540_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n559_), .A2(new_n570_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT71), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n559_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(KEYINPUT13), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  MUX2_X1   g378(.A(new_n245_), .B(new_n247_), .S(new_n292_), .Z(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n292_), .B(new_n245_), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n582_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G113gat), .B(G141gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n583_), .A2(new_n585_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n588_), .B1(new_n592_), .B2(KEYINPUT81), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(KEYINPUT81), .B2(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n579_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n539_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n321_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT101), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n284_), .A3(new_n500_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n278_), .B(KEYINPUT102), .ZN(new_n604_));
  AND4_X1   g403(.A1(new_n319_), .A2(new_n539_), .A3(new_n597_), .A4(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n284_), .B1(new_n605_), .B2(new_n500_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n602_), .B2(new_n601_), .ZN(G1324gat));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n285_), .A3(new_n474_), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT39), .B(new_n285_), .C1(new_n605_), .C2(new_n474_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n474_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n612_), .B2(G8gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g414(.A(new_n605_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n364_), .A2(new_n366_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G15gat), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT103), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(KEYINPUT103), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n620_), .A2(KEYINPUT41), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT41), .B1(new_n620_), .B2(new_n621_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n599_), .A2(G15gat), .A3(new_n617_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT104), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n623_), .A3(new_n625_), .ZN(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n436_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n605_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT42), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n627_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n599_), .B2(new_n631_), .ZN(G1327gat));
  INV_X1    g431(.A(new_n278_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n319_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT106), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(new_n598_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G29gat), .B1(new_n637_), .B2(new_n500_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n535_), .B1(KEYINPUT98), .B2(new_n527_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n628_), .B1(new_n640_), .B2(new_n530_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n617_), .B1(new_n641_), .B2(new_n516_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n281_), .B1(new_n642_), .B2(new_n502_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n639_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n281_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n539_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n597_), .A2(new_n634_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT44), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n653_), .B(new_n650_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n500_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n638_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n636_), .A2(new_n598_), .A3(new_n659_), .A4(new_n474_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT43), .B1(new_n647_), .B2(KEYINPUT105), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n644_), .B(new_n639_), .C1(new_n539_), .C2(new_n646_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n651_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n653_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n474_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n668_), .B2(G36gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n658_), .B1(new_n669_), .B2(KEYINPUT46), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT107), .B(new_n662_), .C1(new_n668_), .C2(G36gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n659_), .B1(new_n655_), .B2(new_n474_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT107), .B1(new_n676_), .B2(new_n662_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n669_), .A2(new_n672_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n677_), .A2(new_n658_), .A3(new_n671_), .A4(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n675_), .A2(new_n679_), .ZN(G1329gat));
  AOI21_X1  g479(.A(G43gat), .B1(new_n637_), .B2(new_n367_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n367_), .A2(G43gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n655_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g483(.A(G50gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n628_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT109), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n637_), .A2(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n652_), .A2(new_n654_), .A3(new_n436_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n685_), .ZN(G1331gat));
  INV_X1    g489(.A(new_n579_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n595_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(new_n539_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n321_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n500_), .ZN(new_n696_));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(KEYINPUT110), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT110), .B1(new_n696_), .B2(new_n697_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n595_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n539_), .A2(new_n604_), .A3(new_n579_), .A4(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n500_), .A2(G57gat), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n699_), .A2(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g504(.A(G64gat), .B1(new_n702_), .B2(new_n475_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT48), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n475_), .A2(G64gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n694_), .B2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n702_), .B2(new_n617_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n617_), .A2(G71gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n694_), .B2(new_n713_), .ZN(G1334gat));
  OAI21_X1  g513(.A(G78gat), .B1(new_n702_), .B2(new_n436_), .ZN(new_n715_));
  XOR2_X1   g514(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n695_), .A2(new_n297_), .A3(new_n628_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1335gat));
  AND3_X1   g518(.A1(new_n649_), .A2(new_n634_), .A3(new_n692_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n202_), .B1(new_n720_), .B2(new_n500_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n693_), .A2(new_n636_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n501_), .A2(G85gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT114), .Z(G1336gat));
  AOI21_X1  g524(.A(new_n203_), .B1(new_n720_), .B2(new_n474_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n475_), .A2(G92gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n722_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT115), .Z(G1337gat));
  AOI21_X1  g528(.A(new_n220_), .B1(new_n720_), .B2(new_n367_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n367_), .A2(new_n209_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n722_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g532(.A1(new_n722_), .A2(new_n210_), .A3(new_n628_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n720_), .A2(new_n628_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G106gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT52), .B(new_n210_), .C1(new_n720_), .C2(new_n628_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g539(.A1(new_n475_), .A2(new_n436_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n617_), .A2(new_n741_), .A3(new_n501_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n581_), .B1(new_n580_), .B2(KEYINPUT118), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(KEYINPUT118), .B2(new_n580_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n588_), .B1(new_n584_), .B2(new_n581_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n591_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n570_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT55), .B1(new_n554_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n565_), .A2(KEYINPUT117), .A3(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n551_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n545_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n545_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(KEYINPUT119), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n760_));
  AOI211_X1 g559(.A(new_n760_), .B(KEYINPUT56), .C1(new_n756_), .C2(new_n545_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n750_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT58), .B(new_n750_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n646_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n595_), .A2(new_n570_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n756_), .A2(new_n545_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n770_), .B2(new_n757_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n748_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n278_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n545_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n595_), .B(new_n570_), .C1(new_n776_), .C2(new_n758_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n772_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT57), .A3(new_n278_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n775_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n634_), .B1(new_n766_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n701_), .A2(new_n578_), .A3(new_n574_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n701_), .A2(new_n574_), .A3(KEYINPUT116), .A4(new_n578_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n281_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT54), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n646_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n743_), .B1(new_n782_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n595_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT120), .Z(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n743_), .B2(KEYINPUT121), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(KEYINPUT121), .B2(new_n743_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT57), .B1(new_n779_), .B2(new_n278_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n774_), .B(new_n633_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n764_), .A2(new_n646_), .A3(new_n765_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n319_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n790_), .B(KEYINPUT54), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n799_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT122), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n806_), .B(KEYINPUT122), .C1(new_n794_), .C2(new_n797_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n596_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n796_), .B1(new_n811_), .B2(new_n813_), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n691_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n794_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n807_), .A2(new_n691_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n819_), .B2(new_n815_), .ZN(G1341gat));
  NAND3_X1  g619(.A1(new_n809_), .A2(new_n319_), .A3(new_n810_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G127gat), .ZN(new_n822_));
  INV_X1    g621(.A(new_n794_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n634_), .A2(G127gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n281_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n809_), .A2(new_n810_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n823_), .B2(new_n604_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT123), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1343gat));
  AOI211_X1 g633(.A(new_n436_), .B(new_n367_), .C1(new_n782_), .C2(new_n793_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(new_n475_), .A3(new_n500_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n596_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n691_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g639(.A1(new_n836_), .A2(new_n634_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT61), .B(G155gat), .Z(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  OAI21_X1  g642(.A(G162gat), .B1(new_n836_), .B2(new_n281_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n604_), .A2(G162gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n836_), .B2(new_n845_), .ZN(G1347gat));
  AOI21_X1  g645(.A(new_n628_), .B1(new_n782_), .B2(new_n793_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n617_), .A2(new_n475_), .A3(new_n500_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n595_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT124), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n851_), .A2(G169gat), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n851_), .B2(G169gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n847_), .A2(new_n848_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n595_), .A2(new_n442_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n853_), .A2(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1348gat));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n691_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n443_), .ZN(G1349gat));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n855_), .A2(new_n634_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n322_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(G183gat), .B2(new_n861_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n860_), .A3(new_n862_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n855_), .B2(new_n281_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n604_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n323_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n855_), .B2(new_n869_), .ZN(G1351gat));
  NAND3_X1  g669(.A1(new_n835_), .A2(new_n474_), .A3(new_n501_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n596_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n370_), .ZN(G1352gat));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n691_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n371_), .ZN(G1353gat));
  NAND2_X1  g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n319_), .A2(new_n876_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT127), .Z(new_n878_));
  NOR2_X1   g677(.A1(new_n871_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1354gat));
  OAI21_X1  g680(.A(G218gat), .B1(new_n871_), .B2(new_n281_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n604_), .A2(G218gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n871_), .B2(new_n883_), .ZN(G1355gat));
endmodule


