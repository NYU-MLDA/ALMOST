//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT90), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G197gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n204_), .A2(new_n205_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n203_), .A2(KEYINPUT90), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(KEYINPUT89), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(KEYINPUT21), .C1(KEYINPUT89), .C2(new_n207_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n203_), .B1(new_n205_), .B2(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n222_), .B2(KEYINPUT1), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n224_), .B2(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT88), .ZN(new_n231_));
  INV_X1    g030(.A(new_n222_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n228_), .B(KEYINPUT3), .Z(new_n233_));
  XOR2_X1   g032(.A(new_n227_), .B(KEYINPUT2), .Z(new_n234_));
  OAI211_X1 g033(.A(new_n220_), .B(new_n232_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n219_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G228gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G78gat), .B(G106gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT91), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n231_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT28), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n231_), .A2(new_n250_), .A3(new_n238_), .A4(new_n235_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n251_), .A3(new_n247_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n245_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n256_), .A2(new_n252_), .A3(new_n242_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n241_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G71gat), .B(G99gat), .ZN(new_n259_));
  INV_X1    g058(.A(G43gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G227gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(G15gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n261_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT24), .A3(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT83), .Z(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT25), .B(G183gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT82), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n268_), .A2(KEYINPUT24), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT23), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n276_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n274_), .A2(KEYINPUT82), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n271_), .A2(new_n275_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n284_), .B(new_n285_), .C1(G183gat), .C2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT22), .B(G169gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT84), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n266_), .A2(KEYINPUT22), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n267_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n286_), .B(new_n269_), .C1(new_n288_), .C2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n283_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n283_), .A2(KEYINPUT30), .A3(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT85), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n299_), .A3(new_n296_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n265_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n265_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G127gat), .B(G134gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n301_), .A2(new_n304_), .A3(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n239_), .B(new_n240_), .Z(new_n315_));
  NAND3_X1  g114(.A1(new_n253_), .A2(new_n243_), .A3(new_n254_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n244_), .B1(new_n256_), .B2(new_n252_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n258_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  OR2_X1    g122(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n236_), .A2(new_n307_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n307_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n231_), .A2(new_n327_), .A3(new_n235_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(KEYINPUT4), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n236_), .A2(new_n330_), .A3(new_n307_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n325_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n325_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n323_), .B(new_n324_), .C1(new_n332_), .C2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n274_), .A2(new_n270_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n338_), .A2(KEYINPUT92), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n281_), .B1(new_n338_), .B2(KEYINPUT92), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n287_), .A2(new_n267_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n286_), .A3(new_n269_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT93), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n212_), .A2(new_n213_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n293_), .A2(new_n219_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(KEYINPUT20), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n219_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n283_), .A3(new_n292_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT20), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n337_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G8gat), .B(G36gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n354_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n323_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n326_), .A2(new_n333_), .A3(new_n328_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n329_), .A2(new_n331_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n361_), .B(new_n362_), .C1(new_n363_), .C2(new_n333_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n335_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n333_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n334_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n324_), .B1(new_n368_), .B2(new_n323_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n346_), .A2(new_n343_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n348_), .B(KEYINPUT20), .C1(new_n341_), .C2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n337_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n350_), .A2(KEYINPUT20), .A3(new_n351_), .A4(new_n373_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n337_), .A2(new_n372_), .B1(new_n374_), .B2(KEYINPUT96), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(KEYINPUT96), .B2(new_n374_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n354_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n377_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n366_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n368_), .A2(new_n323_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n319_), .B1(new_n370_), .B2(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n258_), .A2(new_n318_), .A3(new_n313_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n313_), .B1(new_n258_), .B2(new_n318_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n383_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT97), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n359_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n376_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n380_), .B2(new_n359_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n360_), .A2(KEYINPUT27), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n384_), .A2(KEYINPUT97), .A3(new_n383_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n392_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n386_), .B1(new_n389_), .B2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G29gat), .B(G36gat), .Z(new_n404_));
  XOR2_X1   g203(.A(G43gat), .B(G50gat), .Z(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(KEYINPUT15), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT78), .B(G1gat), .ZN(new_n408_));
  INV_X1    g207(.A(G8gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT14), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G15gat), .B(G22gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G8gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n406_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G229gat), .A2(G233gat), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n418_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n406_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n421_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT81), .Z(new_n426_));
  INV_X1    g225(.A(new_n422_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G113gat), .B(G141gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G169gat), .B(G197gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  OR2_X1    g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n431_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n403_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G190gat), .B(G218gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G134gat), .B(G162gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT36), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G232gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G85gat), .ZN(new_n446_));
  INV_X1    g245(.A(G92gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(KEYINPUT9), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n446_), .A2(new_n447_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n450_), .B(new_n451_), .C1(new_n449_), .C2(KEYINPUT9), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT6), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT10), .B(G99gat), .Z(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n451_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(new_n449_), .A3(KEYINPUT9), .A4(new_n448_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n452_), .A2(new_n454_), .A3(new_n457_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT8), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n454_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n453_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT70), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G99gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n456_), .A3(KEYINPUT67), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(G99gat), .B2(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT68), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n468_), .A2(new_n456_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(KEYINPUT7), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT71), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n469_), .A2(new_n471_), .A3(new_n474_), .A4(new_n472_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n467_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n458_), .A2(new_n448_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT69), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n461_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT68), .B1(new_n486_), .B2(new_n472_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT7), .B1(new_n475_), .B2(new_n470_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(new_n469_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n479_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n454_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n484_), .A2(new_n491_), .A3(new_n461_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n460_), .B(new_n406_), .C1(new_n485_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n460_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n463_), .A2(new_n466_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT71), .B1(new_n489_), .B2(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n484_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT8), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n501_), .B2(new_n492_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n494_), .B1(new_n502_), .B2(new_n407_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n445_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n494_), .B(new_n506_), .C1(new_n502_), .C2(new_n407_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n445_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n441_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n510_), .B2(KEYINPUT76), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT77), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n503_), .A2(new_n504_), .A3(new_n445_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n507_), .B2(new_n505_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n440_), .A2(KEYINPUT36), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(new_n510_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(KEYINPUT37), .C1(new_n510_), .C2(KEYINPUT76), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n517_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526_));
  OR2_X1    g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT79), .Z(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n420_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n531_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT80), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT16), .ZN(new_n538_));
  XOR2_X1   g337(.A(G183gat), .B(G211gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n536_), .A2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n543_), .A2(new_n544_), .B1(new_n534_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n523_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G120gat), .B(G148gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT72), .Z(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n460_), .B1(new_n485_), .B2(new_n493_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n530_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n460_), .B(new_n530_), .C1(new_n485_), .C2(new_n493_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT12), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n555_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n555_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n552_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT73), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n563_), .A2(new_n565_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n551_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NOR4_X1   g369(.A1(new_n563_), .A2(KEYINPUT73), .A3(new_n565_), .A4(new_n551_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT13), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT13), .B(new_n566_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT74), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(KEYINPUT74), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n437_), .A2(new_n547_), .A3(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n392_), .A2(new_n401_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n408_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n432_), .A2(new_n433_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n576_), .A2(new_n546_), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT100), .ZN(new_n588_));
  INV_X1    g387(.A(new_n403_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n517_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(KEYINPUT100), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n588_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n583_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n584_), .A2(new_n585_), .B1(G1gat), .B2(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n584_), .A2(new_n585_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(G1324gat));
  INV_X1    g398(.A(new_n400_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n581_), .A2(new_n409_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n592_), .A2(new_n600_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(G8gat), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT39), .B(new_n409_), .C1(new_n592_), .C2(new_n600_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(G1325gat));
  NAND3_X1  g407(.A1(new_n581_), .A2(new_n263_), .A3(new_n313_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n592_), .A2(new_n313_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n610_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT41), .B1(new_n610_), .B2(G15gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(G1326gat));
  INV_X1    g412(.A(new_n258_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n318_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT102), .Z(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(G22gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT103), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n581_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n592_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G22gat), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT42), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT42), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(G1327gat));
  OR2_X1    g425(.A1(new_n516_), .A2(new_n510_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT76), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n514_), .B2(new_n441_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n518_), .B1(new_n629_), .B2(KEYINPUT37), .ZN(new_n630_));
  INV_X1    g429(.A(new_n519_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n520_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n589_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n523_), .A2(new_n403_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n546_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n576_), .A2(new_n638_), .A3(new_n586_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n639_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(new_n583_), .ZN(new_n645_));
  INV_X1    g444(.A(G29gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n627_), .A2(new_n638_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n576_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n437_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n583_), .A2(new_n646_), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n645_), .A2(new_n646_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  NAND3_X1  g451(.A1(new_n642_), .A2(new_n600_), .A3(new_n643_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n642_), .A2(KEYINPUT104), .A3(new_n600_), .A4(new_n643_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  AND4_X1   g459(.A1(new_n658_), .A2(new_n437_), .A3(new_n600_), .A4(new_n649_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n662_), .B2(new_n661_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n660_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  AOI21_X1  g467(.A(new_n260_), .B1(new_n644_), .B2(new_n313_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n650_), .A2(G43gat), .A3(new_n314_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1330gat));
  INV_X1    g474(.A(G50gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n616_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n437_), .A2(new_n621_), .A3(new_n649_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n644_), .A2(new_n677_), .B1(new_n676_), .B2(new_n678_), .ZN(G1331gat));
  NOR2_X1   g478(.A1(new_n546_), .A2(new_n434_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n590_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n580_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n582_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n403_), .A2(new_n586_), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n685_), .A2(new_n523_), .A3(new_n546_), .A4(new_n577_), .ZN(new_n686_));
  INV_X1    g485(.A(G57gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n583_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n684_), .A2(new_n688_), .ZN(G1332gat));
  OAI21_X1  g488(.A(G64gat), .B1(new_n683_), .B2(new_n400_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n692_), .A3(new_n600_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1333gat));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n695_), .A3(new_n313_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G71gat), .B1(new_n683_), .B2(new_n314_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n699_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(G1334gat));
  INV_X1    g501(.A(G78gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n686_), .A2(new_n703_), .A3(new_n621_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G78gat), .B1(new_n683_), .B2(new_n617_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT50), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT50), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT109), .ZN(G1335gat));
  NOR3_X1   g508(.A1(new_n580_), .A2(new_n648_), .A3(new_n685_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n583_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n577_), .A2(new_n638_), .A3(new_n434_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n637_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n583_), .A2(G85gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT110), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n711_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT111), .ZN(G1336gat));
  AOI21_X1  g517(.A(new_n447_), .B1(new_n714_), .B2(new_n600_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n400_), .A2(G92gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n710_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(G1337gat));
  OAI21_X1  g521(.A(G99gat), .B1(new_n713_), .B2(new_n314_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n313_), .A2(new_n455_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n710_), .A2(new_n724_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n726_), .B(new_n727_), .Z(G1338gat));
  OAI211_X1 g527(.A(new_n710_), .B(new_n456_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  OAI221_X1 g529(.A(G106gat), .B1(KEYINPUT114), .B2(new_n730_), .C1(new_n713_), .C2(new_n616_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT114), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n732_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n729_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  NOR2_X1   g538(.A1(new_n582_), .A2(new_n600_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n387_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n742_));
  INV_X1    g541(.A(new_n570_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n571_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n586_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT116), .B1(new_n563_), .B2(KEYINPUT55), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n559_), .A2(KEYINPUT12), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n501_), .A2(new_n492_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n530_), .B1(new_n748_), .B2(new_n460_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n562_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n564_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n563_), .A2(KEYINPUT55), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n560_), .A2(new_n555_), .A3(new_n562_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n746_), .A2(new_n755_), .A3(new_n756_), .A4(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n758_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT56), .B1(new_n758_), .B2(new_n552_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n745_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n426_), .A2(new_n422_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n431_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n418_), .A2(new_n421_), .A3(new_n427_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n433_), .A2(new_n765_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT117), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n572_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n761_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n742_), .B1(new_n769_), .B2(new_n627_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n771_), .B(new_n517_), .C1(new_n761_), .C2(new_n768_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n743_), .A2(new_n744_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n767_), .B(new_n774_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n776_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n523_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n638_), .B1(new_n773_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n574_), .A2(new_n575_), .A3(new_n680_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n633_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n633_), .B2(new_n782_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n574_), .A2(new_n575_), .A3(new_n680_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n523_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n633_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(KEYINPUT54), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n741_), .B1(new_n780_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(G113gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n434_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT59), .B(new_n741_), .C1(new_n780_), .C2(new_n791_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n586_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n799_), .B2(new_n794_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT119), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n799_), .C2(new_n794_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1340gat));
  INV_X1    g603(.A(G120gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n577_), .B2(KEYINPUT60), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n793_), .B(new_n806_), .C1(KEYINPUT60), .C2(new_n805_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n580_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT120), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n807_), .C1(new_n808_), .C2(new_n805_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1341gat));
  INV_X1    g612(.A(G127gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n793_), .A2(new_n814_), .A3(new_n638_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n546_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n814_), .ZN(G1342gat));
  INV_X1    g616(.A(G134gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n793_), .A2(new_n818_), .A3(new_n517_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n633_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n818_), .ZN(G1343gat));
  INV_X1    g620(.A(new_n388_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n773_), .A2(new_n779_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n546_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n786_), .A2(new_n790_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n822_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n740_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT121), .B1(new_n826_), .B2(new_n740_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n434_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G141gat), .ZN(new_n830_));
  INV_X1    g629(.A(G141gat), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n434_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1344gat));
  OAI21_X1  g632(.A(new_n682_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G148gat), .ZN(new_n835_));
  INV_X1    g634(.A(G148gat), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n682_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1345gat));
  OAI21_X1  g637(.A(new_n638_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n840_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n638_), .B(new_n842_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1346gat));
  INV_X1    g643(.A(G162gat), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n845_), .B(new_n517_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n828_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n740_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n633_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n846_), .B1(new_n849_), .B2(new_n845_), .ZN(G1347gat));
  NAND2_X1  g649(.A1(new_n824_), .A2(new_n825_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n583_), .A2(new_n400_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n313_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n586_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT122), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n617_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G169gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(KEYINPUT62), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n856_), .B2(G169gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n853_), .A2(new_n621_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n851_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n851_), .A2(new_n864_), .A3(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n434_), .A2(new_n287_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n858_), .A2(new_n860_), .B1(new_n866_), .B2(new_n867_), .ZN(G1348gat));
  NAND2_X1  g667(.A1(new_n851_), .A2(new_n616_), .ZN(new_n869_));
  NOR4_X1   g668(.A1(new_n869_), .A2(new_n267_), .A3(new_n580_), .A4(new_n853_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n576_), .A3(new_n865_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n267_), .ZN(G1349gat));
  NOR2_X1   g671(.A1(new_n853_), .A2(new_n546_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n851_), .A2(new_n616_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT124), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(KEYINPUT124), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(G183gat), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n863_), .A2(new_n865_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n546_), .A2(new_n272_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n875_), .A2(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n517_), .A3(new_n273_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G190gat), .B1(new_n866_), .B2(new_n633_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1351gat));
  AND2_X1   g682(.A1(new_n826_), .A2(new_n852_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n434_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n682_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g687(.A(new_n546_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n826_), .A2(new_n852_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n826_), .A2(new_n892_), .A3(new_n852_), .A4(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n895_));
  INV_X1    g694(.A(G211gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n891_), .A2(new_n895_), .A3(new_n896_), .A4(new_n893_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1354gat));
  NAND3_X1  g699(.A1(new_n826_), .A2(new_n517_), .A3(new_n852_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT126), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT127), .B(G218gat), .Z(new_n903_));
  NOR2_X1   g702(.A1(new_n633_), .A2(new_n903_), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n902_), .A2(new_n903_), .B1(new_n884_), .B2(new_n904_), .ZN(G1355gat));
endmodule


