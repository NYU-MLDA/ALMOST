//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT20), .ZN(new_n210_));
  INV_X1    g009(.A(G218gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G211gat), .ZN(new_n212_));
  INV_X1    g011(.A(G211gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G218gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G197gat), .B(G204gat), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n221_));
  INV_X1    g020(.A(G197gat), .ZN(new_n222_));
  INV_X1    g021(.A(G204gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G197gat), .A2(G204gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT91), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n216_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT89), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(KEYINPUT21), .A3(new_n225_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n229_), .B(new_n230_), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT25), .B(G183gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT24), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n235_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT83), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G183gat), .A3(G190gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT23), .ZN(new_n247_));
  OR2_X1    g046(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n248_), .A2(G183gat), .A3(G190gat), .A4(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT23), .B1(new_n244_), .B2(new_n246_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n248_), .A2(new_n249_), .B1(G183gat), .B2(G190gat), .ZN(new_n253_));
  OAI22_X1  g052(.A1(new_n252_), .A2(new_n253_), .B1(G183gat), .B2(G190gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G169gat), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n242_), .A2(new_n251_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n210_), .B1(new_n232_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n235_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n252_), .A2(new_n253_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n256_), .ZN(new_n263_));
  OAI22_X1  g062(.A1(new_n259_), .A2(new_n260_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n209_), .B1(new_n258_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n259_), .A2(new_n260_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n262_), .A2(new_n263_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n218_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n221_), .A2(new_n226_), .A3(KEYINPUT91), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n215_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n229_), .B(new_n230_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n268_), .B(new_n269_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n272_), .A2(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n254_), .A2(new_n256_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n251_), .A2(new_n239_), .A3(new_n241_), .A4(new_n235_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(new_n279_), .A3(KEYINPUT20), .A4(new_n209_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n206_), .B1(new_n267_), .B2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n276_), .B(new_n277_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n265_), .A2(new_n282_), .A3(KEYINPUT20), .A4(new_n209_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT93), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n257_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n275_), .A2(new_n264_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n208_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n258_), .A2(new_n288_), .A3(new_n209_), .A4(new_n265_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n284_), .A2(new_n287_), .A3(new_n289_), .A4(new_n206_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n281_), .B1(KEYINPUT96), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n283_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n274_), .A2(new_n279_), .A3(KEYINPUT20), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n292_), .A2(new_n288_), .B1(new_n293_), .B2(new_n208_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT96), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n206_), .A4(new_n284_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n202_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n284_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n206_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n202_), .A3(new_n290_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT97), .B1(new_n297_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n280_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n299_), .B1(new_n304_), .B2(new_n266_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n290_), .A2(KEYINPUT96), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT27), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT97), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n301_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G22gat), .B(G50gat), .Z(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  INV_X1    g111(.A(G141gat), .ZN(new_n313_));
  INV_X1    g112(.A(G148gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n315_), .A2(new_n318_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  OR2_X1    g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n313_), .A2(new_n314_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n323_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n325_), .B(new_n316_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n324_), .A2(new_n329_), .A3(KEYINPUT86), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT86), .B1(new_n324_), .B2(new_n329_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n311_), .B1(new_n333_), .B2(KEYINPUT29), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  INV_X1    g136(.A(new_n311_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n337_), .B(new_n338_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n324_), .A2(new_n329_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT29), .A3(new_n330_), .ZN(new_n346_));
  INV_X1    g145(.A(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(G228gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(G228gat), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(new_n275_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n343_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n352_), .B1(new_n357_), .B2(new_n232_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G78gat), .B(G106gat), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n363_));
  OAI22_X1  g162(.A1(new_n341_), .A2(new_n342_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n342_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n340_), .A4(new_n361_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT94), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372_));
  XOR2_X1   g171(.A(G127gat), .B(G134gat), .Z(new_n373_));
  XOR2_X1   g172(.A(G113gat), .B(G120gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n345_), .A2(new_n376_), .A3(new_n330_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n355_), .A2(new_n375_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n372_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT4), .B1(new_n333_), .B2(new_n376_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n369_), .B(new_n371_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n331_), .A2(new_n332_), .A3(new_n375_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n376_), .A2(new_n343_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT4), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n377_), .A2(new_n372_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n370_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n377_), .A2(new_n370_), .A3(new_n378_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT94), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n381_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G1gat), .B(G29gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT95), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT0), .B(G57gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n381_), .B(new_n396_), .C1(new_n386_), .C2(new_n388_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT85), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n264_), .B(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n401_), .A2(KEYINPUT31), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(KEYINPUT31), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(G71gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G99gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(new_n375_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n404_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n404_), .A2(new_n411_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n398_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n303_), .A2(new_n310_), .A3(new_n368_), .A4(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n304_), .A2(new_n266_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n418_));
  MUX2_X1   g217(.A(new_n298_), .B(new_n417_), .S(new_n418_), .Z(new_n419_));
  INV_X1    g218(.A(new_n397_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n371_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n388_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n396_), .B1(new_n423_), .B2(new_n381_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n419_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n290_), .B(new_n300_), .C1(new_n424_), .C2(KEYINPUT33), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n389_), .A2(KEYINPUT33), .A3(new_n394_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n370_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n377_), .A2(new_n371_), .A3(new_n378_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n396_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n425_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n308_), .A2(new_n301_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n368_), .A2(new_n398_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n432_), .A2(new_n368_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n414_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n416_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G1gat), .ZN(new_n439_));
  INV_X1    g238(.A(G8gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT77), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT77), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(KEYINPUT14), .C1(new_n439_), .C2(new_n440_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G15gat), .B(G22gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G1gat), .B(G8gat), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n442_), .A2(new_n447_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G29gat), .B(G36gat), .Z(new_n453_));
  XOR2_X1   g252(.A(G43gat), .B(G50gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(KEYINPUT80), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n458_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n452_), .A2(KEYINPUT81), .A3(new_n459_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n459_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(new_n451_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G229gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n451_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n472_));
  INV_X1    g271(.A(new_n458_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n456_), .A2(new_n457_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n455_), .A2(KEYINPUT15), .A3(new_n458_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n463_), .A2(new_n466_), .B1(new_n451_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n471_), .B1(new_n479_), .B2(new_n469_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G169gat), .B(G197gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  OR2_X1    g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G232gat), .A2(G233gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT34), .Z(new_n489_));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G85gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  INV_X1    g301(.A(G99gat), .ZN(new_n503_));
  INV_X1    g302(.A(G106gat), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .A4(KEYINPUT65), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506_));
  OAI22_X1  g305(.A1(new_n506_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n496_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT66), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n507_), .B(new_n505_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n496_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(KEYINPUT8), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n497_), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n504_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n494_), .A2(KEYINPUT9), .A3(new_n495_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n495_), .A2(KEYINPUT9), .ZN(new_n522_));
  AND4_X1   g321(.A1(new_n517_), .A2(new_n520_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n512_), .B1(new_n511_), .B2(new_n496_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n514_), .A2(new_n526_), .A3(new_n460_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n489_), .A2(new_n490_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT71), .Z(new_n529_));
  AOI21_X1  g328(.A(new_n477_), .B1(new_n514_), .B2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n527_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT70), .B(new_n477_), .C1(new_n514_), .C2(new_n526_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n491_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n530_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n491_), .B(KEYINPUT73), .Z(new_n536_));
  NAND4_X1  g335(.A1(new_n535_), .A2(new_n527_), .A3(new_n529_), .A4(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G190gat), .B(G218gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT72), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT37), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n543_), .B(KEYINPUT36), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT74), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n539_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n548_), .B(KEYINPUT74), .Z(new_n552_));
  AND3_X1   g351(.A1(new_n534_), .A2(KEYINPUT75), .A3(new_n537_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT75), .B1(new_n534_), .B2(new_n537_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT76), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT76), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n552_), .B(new_n557_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n546_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n551_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT64), .Z(new_n568_));
  INV_X1    g367(.A(G64gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G57gat), .ZN(new_n570_));
  INV_X1    g369(.A(G57gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(G64gat), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT67), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT11), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n571_), .A2(G64gat), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n569_), .A2(G57gat), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT67), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT11), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G78gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(G71gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n406_), .A2(G78gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n576_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n579_), .A2(new_n581_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(KEYINPUT11), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n514_), .A2(new_n591_), .A3(new_n526_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT68), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n514_), .A2(new_n591_), .A3(new_n526_), .A4(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n514_), .B2(new_n526_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n568_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n568_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n592_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n514_), .A2(new_n526_), .ZN(new_n602_));
  AOI211_X1 g401(.A(new_n580_), .B(new_n586_), .C1(new_n579_), .C2(new_n581_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n589_), .B1(new_n588_), .B2(KEYINPUT11), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n582_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT69), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT12), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n511_), .A2(new_n512_), .A3(new_n496_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n613_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n509_), .A2(KEYINPUT66), .A3(new_n525_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n523_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n605_), .B(new_n612_), .C1(new_n614_), .C2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n601_), .A2(new_n609_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n566_), .B1(new_n598_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n598_), .A2(new_n619_), .A3(new_n566_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT13), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(KEYINPUT13), .A3(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n605_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT78), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n452_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT17), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT17), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n631_), .B(new_n451_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n561_), .A2(new_n628_), .A3(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n438_), .A2(new_n487_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n439_), .A3(new_n398_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n644_), .A2(new_n627_), .A3(new_n487_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n437_), .A2(new_n559_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n398_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n649_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(new_n654_), .A3(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n303_), .A2(new_n310_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n658_), .B(G8gat), .C1(new_n652_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G8gat), .B1(new_n652_), .B2(new_n660_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(KEYINPUT98), .A3(KEYINPUT39), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT98), .B1(new_n664_), .B2(KEYINPUT39), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n663_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n647_), .A2(new_n440_), .A3(new_n659_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n657_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n665_), .A2(new_n666_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT40), .B(new_n668_), .C1(new_n671_), .C2(new_n663_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n647_), .A2(new_n674_), .A3(new_n436_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT100), .ZN(new_n676_));
  INV_X1    g475(.A(new_n652_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n436_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n368_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n647_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n677_), .A2(new_n683_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(G22gat), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n559_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n644_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n627_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n437_), .A3(new_n486_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n398_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n538_), .A2(KEYINPUT36), .A3(new_n544_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT75), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n538_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n534_), .A2(KEYINPUT75), .A3(new_n537_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n549_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n701_), .B2(new_n557_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT37), .B1(new_n702_), .B2(new_n556_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT103), .B1(new_n703_), .B2(new_n551_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n558_), .A2(new_n546_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n699_), .A2(new_n700_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n557_), .B1(new_n706_), .B2(new_n552_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n560_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  INV_X1    g508(.A(new_n551_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n437_), .A2(new_n704_), .A3(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n561_), .A2(KEYINPUT43), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n712_), .A2(KEYINPUT43), .B1(new_n437_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n628_), .A2(new_n486_), .A3(new_n644_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT102), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n696_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n716_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT103), .B(new_n551_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n709_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n719_), .B1(new_n722_), .B2(new_n437_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n713_), .A2(new_n437_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n718_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n717_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n398_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n695_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n717_), .A2(new_n726_), .A3(new_n659_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n693_), .A2(G36gat), .A3(new_n660_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n731_), .A2(KEYINPUT46), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  NAND4_X1  g538(.A1(new_n717_), .A2(new_n726_), .A3(G43gat), .A4(new_n436_), .ZN(new_n740_));
  INV_X1    g539(.A(G43gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n693_), .B2(new_n414_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g543(.A1(new_n717_), .A2(new_n726_), .A3(new_n683_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G50gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n368_), .A2(G50gat), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT105), .Z(new_n748_));
  NAND2_X1  g547(.A1(new_n694_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT106), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n752_), .A3(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n438_), .A2(new_n690_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n628_), .A2(new_n486_), .A3(new_n644_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n757_), .A2(new_n571_), .A3(new_n653_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n438_), .A2(new_n486_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n708_), .A2(new_n710_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(new_n628_), .A3(new_n644_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n763_), .A2(new_n764_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n759_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n767_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT108), .A3(new_n765_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n770_), .A3(new_n398_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n758_), .B1(new_n771_), .B2(new_n571_), .ZN(G1332gat));
  OAI21_X1  g571(.A(G64gat), .B1(new_n757_), .B2(new_n660_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n773_), .A2(KEYINPUT109), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(KEYINPUT109), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n766_), .A2(new_n767_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n569_), .A3(new_n659_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n774_), .A2(KEYINPUT48), .A3(new_n775_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(G1333gat));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n406_), .A3(new_n436_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n755_), .A2(new_n436_), .A3(new_n756_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(G71gat), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G71gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1334gat));
  NAND3_X1  g587(.A1(new_n779_), .A2(new_n583_), .A3(new_n683_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G78gat), .B1(new_n757_), .B2(new_n368_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT50), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(KEYINPUT50), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(G1335gat));
  NAND3_X1  g592(.A1(new_n644_), .A2(new_n627_), .A3(new_n487_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n714_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n653_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n438_), .A2(new_n486_), .A3(new_n628_), .A4(new_n691_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n492_), .A3(new_n398_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1336gat));
  OAI21_X1  g599(.A(G92gat), .B1(new_n796_), .B2(new_n660_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n493_), .A3(new_n659_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1337gat));
  NAND4_X1  g602(.A1(new_n798_), .A2(new_n436_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n794_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n436_), .B(new_n805_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT111), .B1(new_n806_), .B2(G99gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT51), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n804_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n798_), .A2(new_n504_), .A3(new_n683_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n683_), .B(new_n805_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(G106gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT53), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n814_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1339gat));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n467_), .A2(new_n470_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n483_), .B1(new_n825_), .B2(new_n468_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n479_), .A2(new_n469_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n480_), .A2(new_n483_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n623_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n622_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n828_), .B(new_n824_), .C1(new_n830_), .C2(new_n620_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n618_), .B1(new_n597_), .B2(new_n607_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n568_), .B1(new_n834_), .B2(new_n596_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n834_), .B2(new_n600_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n601_), .A2(new_n609_), .A3(KEYINPUT55), .A4(new_n618_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n565_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT112), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n843_), .A3(new_n565_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n841_), .A2(KEYINPUT113), .A3(new_n842_), .A4(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n830_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n839_), .A2(KEYINPUT56), .A3(new_n565_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n843_), .B1(new_n839_), .B2(new_n565_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(KEYINPUT56), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n844_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n833_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT57), .A3(new_n559_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n848_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n839_), .B2(new_n565_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n622_), .B(new_n828_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n859_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n761_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n844_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n863_), .A2(new_n851_), .A3(KEYINPUT56), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n845_), .B(new_n846_), .C1(new_n864_), .C2(new_n850_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n690_), .B1(new_n865_), .B2(new_n833_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n867_));
  OAI211_X1 g666(.A(new_n855_), .B(new_n862_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n646_), .B2(new_n486_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n703_), .A2(new_n644_), .A3(new_n551_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n487_), .A4(new_n628_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n868_), .A2(new_n644_), .B1(new_n869_), .B2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n659_), .A2(new_n683_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n436_), .A3(new_n398_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n486_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n873_), .B2(new_n875_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n875_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n858_), .B(KEYINPUT58), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n866_), .A2(KEYINPUT57), .B1(new_n882_), .B2(new_n761_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n854_), .A2(new_n559_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n867_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n645_), .B1(new_n883_), .B2(new_n886_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n869_), .A2(new_n872_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n880_), .B(new_n881_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n879_), .A2(KEYINPUT117), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n876_), .A2(new_n891_), .A3(new_n881_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n487_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n878_), .B1(new_n893_), .B2(new_n877_), .ZN(G1340gat));
  NAND2_X1  g693(.A1(new_n868_), .A2(new_n644_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n869_), .A2(new_n872_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898_));
  AOI21_X1  g697(.A(G120gat), .B1(new_n627_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n898_), .B2(G120gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(new_n880_), .A3(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT118), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n628_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n903_));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n876_), .A2(new_n906_), .A3(new_n645_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n644_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(G1342gat));
  INV_X1    g708(.A(G134gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n876_), .A2(new_n910_), .A3(new_n690_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n561_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(G1343gat));
  NOR2_X1   g712(.A1(new_n436_), .A2(new_n368_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR4_X1   g714(.A1(new_n873_), .A2(new_n653_), .A3(new_n659_), .A4(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n486_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n627_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT119), .B(G148gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1345gat));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n645_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  AOI21_X1  g723(.A(G162gat), .B1(new_n916_), .B2(new_n690_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n722_), .A2(G162gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n916_), .B2(new_n926_), .ZN(G1347gat));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n659_), .A2(new_n368_), .A3(new_n415_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n897_), .A2(new_n486_), .A3(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  AND4_X1   g730(.A1(new_n928_), .A2(new_n930_), .A3(new_n931_), .A4(G169gat), .ZN(new_n932_));
  INV_X1    g731(.A(G169gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(KEYINPUT120), .B2(KEYINPUT62), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n930_), .A2(new_n934_), .B1(new_n928_), .B2(new_n931_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT22), .B(G169gat), .Z(new_n936_));
  OAI22_X1  g735(.A1(new_n932_), .A2(new_n935_), .B1(new_n930_), .B2(new_n936_), .ZN(G1348gat));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938_));
  INV_X1    g737(.A(G176gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n628_), .B1(KEYINPUT121), .B2(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n929_), .B(new_n940_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT122), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n897_), .A2(new_n943_), .A3(new_n929_), .A4(new_n940_), .ZN(new_n944_));
  AND4_X1   g743(.A1(new_n938_), .A2(new_n942_), .A3(new_n944_), .A4(G176gat), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n942_), .A2(new_n944_), .B1(new_n938_), .B2(G176gat), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1349gat));
  NAND2_X1  g746(.A1(new_n897_), .A2(new_n929_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n644_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n949_), .B(new_n233_), .C1(KEYINPUT123), .C2(G183gat), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(G183gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n950_), .B1(new_n949_), .B2(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n948_), .B2(new_n561_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n690_), .A2(new_n234_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n948_), .B2(new_n955_), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n660_), .A2(new_n398_), .A3(new_n915_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(KEYINPUT124), .B1(new_n873_), .B2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n960_), .B(new_n957_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n222_), .A2(KEYINPUT125), .ZN(new_n963_));
  AND3_X1   g762(.A1(new_n962_), .A2(new_n486_), .A3(new_n963_), .ZN(new_n964_));
  OR2_X1    g763(.A1(new_n222_), .A2(KEYINPUT125), .ZN(new_n965_));
  AOI22_X1  g764(.A1(new_n962_), .A2(new_n486_), .B1(new_n965_), .B2(new_n963_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1352gat));
  AOI21_X1  g766(.A(new_n628_), .B1(new_n959_), .B2(new_n961_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(new_n223_), .ZN(G1353gat));
  AOI21_X1  g768(.A(new_n644_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n970_));
  OR3_X1    g769(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971_));
  AND3_X1   g770(.A1(new_n962_), .A2(new_n970_), .A3(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  AOI22_X1  g772(.A1(new_n962_), .A2(new_n970_), .B1(new_n973_), .B2(new_n971_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n972_), .A2(new_n974_), .ZN(G1354gat));
  NAND3_X1  g774(.A1(new_n962_), .A2(new_n211_), .A3(new_n690_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n561_), .B1(new_n959_), .B2(new_n961_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n211_), .ZN(G1355gat));
endmodule


