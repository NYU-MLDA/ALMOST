//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n826_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT66), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n216_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(KEYINPUT67), .A3(new_n216_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT8), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT8), .B1(new_n211_), .B2(new_n212_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n208_), .A2(new_n209_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n225_), .A2(KEYINPUT65), .A3(new_n210_), .A4(new_n205_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .A4(new_n216_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G50gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT69), .B(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT10), .B(G99gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n204_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT9), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .A4(new_n225_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n229_), .A2(new_n233_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT34), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT35), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n244_), .A2(new_n245_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n233_), .B(KEYINPUT15), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n229_), .A2(new_n240_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT73), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n247_), .A2(KEYINPUT70), .B1(new_n250_), .B2(new_n251_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(KEYINPUT70), .B2(new_n247_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n248_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G190gat), .B(G218gat), .ZN(new_n259_));
  INV_X1    g058(.A(G162gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT71), .B(G134gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n265_), .B(KEYINPUT72), .Z(new_n268_));
  NAND3_X1  g067(.A1(new_n254_), .A2(new_n257_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT74), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n269_), .A2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n267_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G15gat), .B(G22gat), .Z(new_n276_));
  NAND2_X1  g075(.A1(G1gat), .A2(G8gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n276_), .B1(KEYINPUT14), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT75), .ZN(new_n279_));
  XOR2_X1   g078(.A(G1gat), .B(G8gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n278_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G231gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G78gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n294_), .B2(new_n291_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n288_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G127gat), .B(G155gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G211gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT16), .B(G183gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n303_));
  OR3_X1    g102(.A1(new_n297_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n302_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(KEYINPUT76), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n306_), .B1(KEYINPUT76), .B2(new_n304_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n275_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT77), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n315_), .A2(KEYINPUT24), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT23), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n318_), .B(new_n320_), .C1(KEYINPUT24), .C2(new_n313_), .ZN(new_n321_));
  OR2_X1    g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n320_), .A2(new_n322_), .B1(G169gat), .B2(G176gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT83), .B1(new_n324_), .B2(G169gat), .ZN(new_n325_));
  INV_X1    g124(.A(G176gat), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n324_), .A2(G169gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(G169gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n326_), .B(new_n327_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n323_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n321_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G15gat), .B(G43gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT84), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT31), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT30), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n340_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n334_), .B(new_n344_), .Z(new_n345_));
  XOR2_X1   g144(.A(G141gat), .B(G148gat), .Z(new_n346_));
  INV_X1    g145(.A(G155gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT1), .B1(new_n347_), .B2(new_n260_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(G155gat), .B2(G162gat), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n347_), .A2(new_n260_), .A3(KEYINPUT1), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n346_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n347_), .A2(new_n260_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359_));
  OAI22_X1  g158(.A1(new_n356_), .A2(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n358_), .B(new_n359_), .C1(G141gat), .C2(G148gat), .ZN(new_n361_));
  INV_X1    g160(.A(G141gat), .ZN(new_n362_));
  INV_X1    g161(.A(G148gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n363_), .C1(KEYINPUT86), .C2(KEYINPUT3), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n356_), .A2(new_n357_), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n354_), .B(new_n355_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n353_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n339_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT4), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n368_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G85gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(new_n238_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT18), .B(G64gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G204gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(G197gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT87), .B(G197gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n393_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT21), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT88), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G197gat), .A2(G204gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT21), .B(new_n401_), .C1(new_n395_), .C2(G204gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(KEYINPUT21), .A3(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n332_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n311_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n318_), .B(new_n320_), .C1(KEYINPUT24), .C2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n327_), .A2(new_n328_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n323_), .B1(G176gat), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT20), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n414_), .B2(KEYINPUT90), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n416_), .A3(KEYINPUT20), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n392_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n412_), .A2(new_n405_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(KEYINPUT20), .C1(new_n332_), .C2(new_n405_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n391_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n389_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n406_), .A2(new_n391_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(KEYINPUT20), .A3(new_n413_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n389_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n391_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(KEYINPUT27), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n405_), .B1(new_n368_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n431_), .B(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G78gat), .B(G106gat), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT89), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n368_), .A2(new_n430_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G22gat), .B(G50gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT28), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n439_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n434_), .A2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n437_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n438_), .A2(new_n444_), .A3(new_n437_), .A4(new_n442_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n425_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n427_), .B2(new_n450_), .ZN(new_n451_));
  AND4_X1   g250(.A1(new_n385_), .A2(new_n429_), .A3(new_n448_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n424_), .A2(new_n453_), .A3(new_n426_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n455_), .B(new_n456_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n383_), .A2(KEYINPUT33), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n427_), .A2(new_n450_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n370_), .A2(new_n373_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n382_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n448_), .B1(new_n457_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n345_), .B1(new_n452_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n429_), .A2(new_n451_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(new_n448_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n385_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n345_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n310_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n286_), .A2(new_n233_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n283_), .A2(new_n284_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n279_), .A2(new_n280_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n233_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT78), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n286_), .A2(KEYINPUT78), .A3(new_n233_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n475_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT79), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n286_), .A2(KEYINPUT78), .A3(new_n233_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT78), .B1(new_n286_), .B2(new_n233_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n485_), .A2(new_n486_), .B1(new_n233_), .B2(new_n286_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488_));
  INV_X1    g287(.A(new_n483_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n484_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n250_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(new_n483_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT80), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n480_), .A2(new_n481_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n483_), .A4(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT81), .B(G169gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G197gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n251_), .A2(new_n295_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT12), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT68), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n229_), .A2(new_n240_), .A3(new_n296_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(KEYINPUT68), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT64), .Z(new_n518_));
  NAND3_X1  g317(.A1(new_n251_), .A2(new_n295_), .A3(new_n511_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n513_), .A2(new_n516_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n509_), .A2(new_n514_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT5), .B(G176gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n393_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G120gat), .B(G148gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n522_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n522_), .A2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n526_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT13), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n508_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n474_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G1gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n470_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT38), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT93), .Z(new_n541_));
  NAND3_X1  g340(.A1(new_n473_), .A2(new_n307_), .A3(new_n273_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n535_), .B(KEYINPUT92), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n537_), .B1(new_n545_), .B2(new_n470_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n538_), .A2(new_n547_), .A3(new_n539_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n550_), .ZN(G1324gat));
  INV_X1    g350(.A(G8gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n545_), .B2(new_n468_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT39), .Z(new_n554_));
  NAND3_X1  g353(.A1(new_n536_), .A2(new_n552_), .A3(new_n468_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT94), .B(KEYINPUT40), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(G1325gat));
  INV_X1    g357(.A(G15gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n345_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n545_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT41), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n536_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(G1326gat));
  INV_X1    g363(.A(G22gat), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n545_), .B2(new_n448_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT42), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n536_), .A2(new_n565_), .A3(new_n448_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT95), .Z(G1327gat));
  INV_X1    g369(.A(G29gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n544_), .A2(new_n308_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT96), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n544_), .A2(new_n574_), .A3(new_n308_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT43), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n473_), .A2(new_n576_), .A3(new_n275_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n473_), .B2(new_n275_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n573_), .B(new_n575_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT97), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT44), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(KEYINPUT97), .A3(KEYINPUT44), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n571_), .B1(new_n585_), .B2(new_n470_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT98), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n273_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n308_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(new_n508_), .A3(new_n534_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n571_), .A3(new_n470_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(G1328gat));
  INV_X1    g391(.A(G36gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n593_), .A3(new_n468_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n585_), .A2(new_n468_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(G36gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(KEYINPUT46), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n598_), .A2(KEYINPUT101), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n594_), .B(new_n595_), .Z(new_n602_));
  INV_X1    g401(.A(new_n468_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n604_), .B2(new_n593_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n599_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n602_), .B(KEYINPUT46), .C1(new_n604_), .C2(new_n593_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(KEYINPUT102), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(KEYINPUT102), .ZN(new_n610_));
  OAI22_X1  g409(.A1(new_n600_), .A2(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(G1329gat));
  INV_X1    g410(.A(new_n590_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n612_), .A2(G43gat), .A3(new_n345_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n585_), .A2(new_n560_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n614_), .B2(G43gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g415(.A(G50gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n590_), .A2(new_n617_), .A3(new_n448_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n448_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n620_), .B2(new_n617_), .ZN(G1331gat));
  AND2_X1   g420(.A1(new_n529_), .A2(new_n533_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n507_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n543_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT104), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(G57gat), .A3(new_n470_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n474_), .A2(new_n623_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G57gat), .B1(new_n627_), .B2(new_n470_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(G1332gat));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n468_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(G64gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n633_), .B2(G64gat), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT48), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT106), .B1(new_n603_), .B2(G64gat), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n603_), .A2(KEYINPUT106), .A3(G64gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n641_), .A3(new_n642_), .ZN(G1333gat));
  INV_X1    g442(.A(G71gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n625_), .B2(new_n560_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT49), .Z(new_n646_));
  NOR2_X1   g445(.A1(new_n345_), .A2(G71gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT107), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n627_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1334gat));
  INV_X1    g449(.A(G78gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n625_), .B2(new_n448_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT50), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n627_), .A2(new_n651_), .A3(new_n448_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1335gat));
  OAI211_X1 g454(.A(new_n308_), .B(new_n623_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT109), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(G85gat), .A3(new_n470_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n588_), .A2(new_n308_), .A3(new_n623_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT108), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n237_), .B1(new_n660_), .B2(new_n385_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n658_), .A2(new_n661_), .ZN(G1336gat));
  INV_X1    g461(.A(new_n660_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G92gat), .B1(new_n663_), .B2(new_n468_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n603_), .A2(new_n238_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n657_), .B2(new_n665_), .ZN(G1337gat));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n234_), .A3(new_n560_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n657_), .A2(new_n560_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(new_n203_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g469(.A(G106gat), .B1(new_n656_), .B2(new_n619_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT52), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n204_), .A3(new_n448_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g474(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n676_));
  NAND2_X1  g475(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n307_), .A2(new_n622_), .A3(new_n508_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT110), .Z(new_n680_));
  INV_X1    g479(.A(new_n275_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n676_), .B(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n680_), .A2(new_n681_), .A3(new_n678_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n492_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT117), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT117), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n495_), .A2(new_n687_), .A3(new_n492_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n489_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n487_), .A2(new_n483_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n504_), .A3(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n506_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n511_), .B1(new_n251_), .B2(new_n295_), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n296_), .B(new_n512_), .C1(new_n229_), .C2(new_n240_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n518_), .B1(new_n695_), .B2(new_n516_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n520_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n698_), .B2(KEYINPUT113), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n520_), .A2(new_n700_), .A3(new_n697_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT55), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT114), .B1(new_n520_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n514_), .A2(new_n515_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n693_), .A2(new_n694_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT114), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(KEYINPUT55), .A4(new_n518_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n699_), .A2(new_n701_), .A3(new_n703_), .A4(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT56), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n526_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n692_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n708_), .B2(new_n526_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n530_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT58), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT120), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT120), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n711_), .A2(new_n713_), .A3(new_n719_), .A4(KEYINPUT58), .ZN(new_n720_));
  AND4_X1   g519(.A1(new_n275_), .A2(new_n716_), .A3(new_n718_), .A4(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n698_), .A2(KEYINPUT113), .ZN(new_n722_));
  INV_X1    g521(.A(new_n696_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(new_n703_), .A3(new_n707_), .A4(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n701_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n526_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n531_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT115), .B1(new_n708_), .B2(new_n526_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n507_), .B1(new_n730_), .B2(KEYINPUT56), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT116), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n530_), .B1(new_n712_), .B2(new_n727_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n726_), .A2(new_n727_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n709_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n733_), .A2(new_n735_), .A3(new_n736_), .A4(new_n507_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n692_), .A2(KEYINPUT118), .A3(new_n527_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT118), .B1(new_n692_), .B2(new_n527_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n732_), .A2(new_n737_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n273_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n741_), .A2(new_n744_), .A3(new_n273_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n721_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n308_), .B1(new_n746_), .B2(KEYINPUT121), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n275_), .A2(new_n716_), .A3(new_n718_), .A4(new_n720_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n741_), .A2(new_n744_), .A3(new_n273_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n741_), .B2(new_n273_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT121), .B(new_n748_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n684_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n469_), .A2(new_n470_), .A3(new_n560_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT122), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT59), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n308_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n684_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n755_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n757_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(G113gat), .A3(new_n507_), .ZN(new_n764_));
  INV_X1    g563(.A(G113gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n756_), .B2(new_n508_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1340gat));
  INV_X1    g566(.A(G120gat), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT60), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n753_), .A2(new_n755_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT123), .ZN(new_n772_));
  INV_X1    g571(.A(new_n755_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n758_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n308_), .A3(new_n751_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n773_), .B1(new_n776_), .B2(new_n684_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT123), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n534_), .B(new_n762_), .C1(new_n777_), .C2(new_n761_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G120gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT124), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n782_), .A3(KEYINPUT124), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1341gat));
  NAND3_X1  g586(.A1(new_n763_), .A2(G127gat), .A3(new_n307_), .ZN(new_n788_));
  INV_X1    g587(.A(G127gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n756_), .B2(new_n308_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1342gat));
  NAND3_X1  g590(.A1(new_n763_), .A2(G134gat), .A3(new_n275_), .ZN(new_n792_));
  INV_X1    g591(.A(G134gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n756_), .B2(new_n273_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1343gat));
  NOR2_X1   g594(.A1(new_n468_), .A2(new_n619_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n753_), .A2(new_n470_), .A3(new_n345_), .A4(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n508_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(new_n362_), .ZN(G1344gat));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n622_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(new_n363_), .ZN(G1345gat));
  XNOR2_X1  g600(.A(KEYINPUT61), .B(G155gat), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT125), .B1(new_n797_), .B2(new_n308_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n797_), .A2(KEYINPUT125), .A3(new_n308_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n804_), .A3(new_n802_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1346gat));
  NOR3_X1   g609(.A1(new_n797_), .A2(new_n260_), .A3(new_n681_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n797_), .A2(new_n273_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n260_), .B2(new_n812_), .ZN(G1347gat));
  NAND3_X1  g612(.A1(new_n471_), .A2(new_n468_), .A3(new_n619_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n684_), .B2(new_n759_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G169gat), .B1(new_n816_), .B2(new_n508_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n507_), .A3(new_n409_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n818_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(G1348gat));
  NAND3_X1  g621(.A1(new_n815_), .A2(new_n326_), .A3(new_n534_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n622_), .B(new_n814_), .C1(new_n776_), .C2(new_n684_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n326_), .ZN(G1349gat));
  NAND2_X1  g624(.A1(new_n815_), .A2(new_n307_), .ZN(new_n826_));
  MUX2_X1   g625(.A(new_n316_), .B(G183gat), .S(new_n826_), .Z(G1350gat));
  OAI21_X1  g626(.A(G190gat), .B1(new_n816_), .B2(new_n681_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n273_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n317_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n816_), .B2(new_n830_), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT126), .Z(G1351gat));
  AOI21_X1  g631(.A(new_n560_), .B1(new_n776_), .B2(new_n684_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n603_), .A2(new_n470_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n448_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n507_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n833_), .A2(new_n507_), .A3(new_n448_), .A4(new_n834_), .ZN(new_n838_));
  INV_X1    g637(.A(G197gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT127), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n837_), .A2(new_n840_), .A3(new_n842_), .ZN(G1352gat));
  NOR2_X1   g642(.A1(new_n835_), .A2(new_n622_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n393_), .ZN(G1353gat));
  NOR2_X1   g644(.A1(new_n835_), .A2(new_n308_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n847_));
  AND2_X1   g646(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n846_), .B2(new_n847_), .ZN(G1354gat));
  AOI21_X1  g649(.A(G218gat), .B1(new_n836_), .B2(new_n829_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n835_), .A2(new_n681_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(G218gat), .B2(new_n852_), .ZN(G1355gat));
endmodule


