//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT25), .B(G183gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n209_), .A2(KEYINPUT79), .A3(new_n212_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT23), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n204_), .B2(KEYINPUT24), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(KEYINPUT80), .B(new_n218_), .C1(new_n204_), .C2(KEYINPUT24), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n215_), .A2(new_n216_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT81), .B(G176gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n208_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G99gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G43gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n229_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n232_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n237_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT82), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G155gat), .A3(G162gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G155gat), .ZN(new_n254_));
  INV_X1    g053(.A(G162gat), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n253_), .A2(KEYINPUT1), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(KEYINPUT1), .B2(new_n253_), .ZN(new_n257_));
  AND2_X1   g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(KEYINPUT83), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n258_), .A2(KEYINPUT2), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n258_), .A2(KEYINPUT2), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n250_), .A2(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n265_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT29), .ZN(new_n275_));
  INV_X1    g074(.A(G197gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G204gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT86), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n280_));
  INV_X1    g079(.A(G204gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G197gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT85), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n279_), .A2(new_n280_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G211gat), .B(G218gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n277_), .A2(new_n282_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(KEYINPUT21), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n279_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT88), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n286_), .A2(new_n289_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT88), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(G228gat), .A2(G233gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n248_), .B1(new_n275_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n275_), .A2(new_n301_), .A3(new_n248_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n275_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n300_), .B1(new_n306_), .B2(new_n296_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G78gat), .B(G106gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n263_), .A2(new_n264_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G22gat), .B(G50gat), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n313_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n309_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n305_), .A2(new_n319_), .A3(new_n307_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n310_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n318_), .B1(new_n310_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n247_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n236_), .B1(new_n274_), .B2(KEYINPUT98), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT98), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n311_), .A2(new_n326_), .A3(new_n235_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT4), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n274_), .A2(new_n330_), .A3(new_n235_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(KEYINPUT99), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n330_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(new_n334_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G85gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT0), .B(G57gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n328_), .A2(new_n332_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n336_), .A2(new_n339_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT100), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n336_), .A2(new_n344_), .A3(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n346_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n226_), .B(KEYINPUT93), .Z(new_n357_));
  AOI22_X1  g156(.A1(new_n357_), .A2(new_n225_), .B1(new_n224_), .B2(KEYINPUT94), .ZN(new_n358_));
  INV_X1    g157(.A(new_n224_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n207_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n208_), .B2(new_n203_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT92), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n218_), .A3(new_n212_), .A4(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n296_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT20), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n295_), .A2(new_n298_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n229_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT95), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n229_), .A2(KEYINPUT95), .A3(new_n295_), .A4(new_n298_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n356_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n362_), .A2(new_n369_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n294_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n379_), .B(KEYINPUT20), .C1(new_n372_), .C2(new_n229_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n355_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n375_), .A2(KEYINPUT96), .A3(new_n356_), .A4(new_n376_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n228_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n209_), .A2(KEYINPUT79), .A3(new_n212_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT79), .B1(new_n209_), .B2(new_n212_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n221_), .A2(new_n222_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n374_), .B1(new_n299_), .B2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n370_), .A2(KEYINPUT20), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n356_), .A4(new_n376_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(new_n355_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n383_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n402_));
  MUX2_X1   g201(.A(new_n382_), .B(new_n396_), .S(new_n402_), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n352_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n345_), .B(KEYINPUT33), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n392_), .A2(new_n393_), .B1(new_n355_), .B2(new_n380_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n406_), .A2(new_n401_), .A3(new_n383_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n401_), .B1(new_n406_), .B2(new_n383_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n343_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n331_), .A2(new_n332_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n338_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n324_), .B1(new_n404_), .B2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n316_), .B(new_n317_), .Z(new_n415_));
  AND3_X1   g214(.A1(new_n305_), .A2(new_n319_), .A3(new_n307_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n319_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n247_), .B1(new_n418_), .B2(new_n321_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n401_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n396_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n406_), .A2(new_n401_), .A3(new_n383_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT27), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n420_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT27), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT101), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT27), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT101), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n419_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n418_), .A2(new_n321_), .A3(new_n247_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n423_), .A2(new_n425_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n352_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n414_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G22gat), .ZN(new_n440_));
  INV_X1    g239(.A(G1gat), .ZN(new_n441_));
  INV_X1    g240(.A(G8gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT14), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G8gat), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449_));
  INV_X1    g248(.A(G29gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(G36gat), .ZN(new_n451_));
  INV_X1    g250(.A(G36gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(G29gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(G29gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(G36gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT68), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G43gat), .B(G50gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n448_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n448_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT76), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT76), .ZN(new_n466_));
  INV_X1    g265(.A(new_n464_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n462_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n454_), .A2(new_n457_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n458_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n459_), .A3(KEYINPUT15), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n448_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n462_), .A2(new_n471_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n469_), .A2(new_n471_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT77), .ZN(new_n483_));
  XOR2_X1   g282(.A(G169gat), .B(G197gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n481_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n439_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G190gat), .B(G218gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT71), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G134gat), .B(G162gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT36), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n494_), .B(KEYINPUT73), .Z(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  INV_X1    g300(.A(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(KEYINPUT9), .ZN(new_n506_));
  INV_X1    g305(.A(G85gat), .ZN(new_n507_));
  INV_X1    g306(.A(G92gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT9), .A3(new_n505_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n500_), .A2(new_n504_), .A3(new_n506_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n502_), .A4(KEYINPUT64), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n515_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n514_), .A2(new_n516_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT8), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n509_), .A2(new_n505_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n511_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT65), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n460_), .A2(new_n461_), .ZN(new_n525_));
  OAI211_X1 g324(.A(KEYINPUT65), .B(new_n511_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n478_), .A2(new_n522_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n527_), .A2(new_n533_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n527_), .A2(new_n534_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT69), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n527_), .A2(KEYINPUT69), .A3(new_n534_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n533_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AOI211_X1 g345(.A(KEYINPUT70), .B(new_n533_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n495_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n541_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n543_), .A3(new_n535_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n532_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT70), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n544_), .A2(new_n545_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n493_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .A4(new_n538_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n489_), .B1(new_n548_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT74), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n548_), .B2(new_n557_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  OAI22_X1  g360(.A1(KEYINPUT74), .A2(new_n558_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n495_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n536_), .B(KEYINPUT72), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n551_), .B2(KEYINPUT70), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n565_), .B2(new_n553_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n546_), .A2(new_n555_), .A3(new_n547_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT75), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n559_), .A3(KEYINPUT37), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G78gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G78gat), .B1(new_n577_), .B2(new_n572_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(G57gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(G64gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n580_), .A2(G64gat), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(KEYINPUT11), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT11), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n583_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n581_), .A3(KEYINPUT11), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n587_), .A2(new_n589_), .A3(new_n578_), .A4(new_n576_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n517_), .A2(new_n519_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT8), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT65), .B1(new_n596_), .B2(new_n511_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n526_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n592_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n524_), .A2(new_n526_), .A3(new_n591_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n511_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n585_), .A2(new_n590_), .A3(KEYINPUT12), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT67), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n585_), .A2(new_n590_), .A3(KEYINPUT12), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT67), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n522_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n591_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n612_), .B(new_n600_), .C1(new_n613_), .C2(KEYINPUT12), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n604_), .B1(new_n614_), .B2(new_n603_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n604_), .B(new_n621_), .C1(new_n614_), .C2(new_n603_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT13), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n623_), .A2(new_n624_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n591_), .B(new_n448_), .Z(new_n630_));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT16), .ZN(new_n634_));
  XOR2_X1   g433(.A(G183gat), .B(G211gat), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT17), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n632_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT17), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n641_), .B2(new_n632_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n571_), .A2(new_n629_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n488_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n352_), .A2(new_n441_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n404_), .A2(new_n413_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n324_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n426_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n429_), .A2(KEYINPUT101), .A3(new_n430_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n655_), .A2(new_n419_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n656_), .B2(new_n352_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n628_), .A2(new_n486_), .A3(new_n642_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT102), .Z(new_n659_));
  NOR2_X1   g458(.A1(new_n566_), .A2(new_n567_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n438_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n649_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT103), .ZN(G1324gat));
  INV_X1    g463(.A(new_n660_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n439_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n655_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(KEYINPUT105), .A3(new_n667_), .A4(new_n659_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n661_), .B2(new_n655_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n670_), .A3(G8gat), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n655_), .A2(G8gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n488_), .A2(new_n644_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n488_), .A2(new_n676_), .A3(new_n644_), .A4(new_n673_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n671_), .A2(new_n672_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n668_), .A2(new_n670_), .A3(KEYINPUT39), .A4(G8gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n247_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n666_), .A2(new_n684_), .A3(new_n659_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT41), .B1(new_n685_), .B2(G15gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n240_), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n686_), .A2(new_n687_), .B1(new_n645_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n322_), .A2(new_n323_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G22gat), .B1(new_n661_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT42), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n693_), .A2(G22gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n645_), .B2(new_n696_), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n665_), .A2(new_n643_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n629_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n488_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n450_), .B1(new_n700_), .B2(new_n438_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n629_), .A2(new_n487_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n643_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n570_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n657_), .A2(new_n705_), .A3(new_n571_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(G29gat), .B(new_n352_), .C1(new_n707_), .C2(KEYINPUT44), .ZN(new_n708_));
  INV_X1    g507(.A(new_n703_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n439_), .A2(KEYINPUT43), .A3(new_n570_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n705_), .B1(new_n657_), .B2(new_n571_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n701_), .B1(new_n708_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT108), .ZN(G1328gat));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n667_), .A2(new_n452_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n700_), .A2(KEYINPUT45), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT45), .B1(new_n700_), .B2(new_n718_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n655_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n707_), .A2(KEYINPUT44), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n452_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n717_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n667_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n727_));
  OAI21_X1  g526(.A(G36gat), .B1(new_n727_), .B2(new_n714_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(KEYINPUT46), .A3(new_n721_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1329gat));
  OAI211_X1 g529(.A(G43gat), .B(new_n684_), .C1(new_n707_), .C2(KEYINPUT44), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n700_), .A2(new_n247_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n731_), .A2(new_n714_), .B1(G43gat), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g533(.A1(new_n700_), .A2(G50gat), .A3(new_n693_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n692_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n714_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G50gat), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n737_), .A2(new_n714_), .A3(new_n736_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(G1331gat));
  NOR2_X1   g540(.A1(new_n643_), .A2(new_n486_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n666_), .A2(new_n629_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n438_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n439_), .A2(new_n486_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n570_), .A2(new_n629_), .A3(new_n642_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n352_), .A2(new_n580_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n743_), .B2(new_n655_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT48), .Z(new_n754_));
  NOR3_X1   g553(.A1(new_n750_), .A2(G64gat), .A3(new_n655_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n743_), .B2(new_n247_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n247_), .A2(G71gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT111), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n750_), .B2(new_n760_), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n743_), .B2(new_n693_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n692_), .A2(new_n574_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n763_), .A2(new_n764_), .B1(new_n750_), .B2(new_n765_), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n698_), .A2(new_n628_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n745_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n507_), .A3(new_n352_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n628_), .A2(new_n486_), .A3(new_n642_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(new_n352_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n774_), .B2(new_n507_), .ZN(G1336gat));
  NAND3_X1  g574(.A1(new_n769_), .A2(new_n508_), .A3(new_n667_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n773_), .A2(new_n667_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n508_), .ZN(G1337gat));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n501_), .A2(new_n503_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n684_), .A2(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n745_), .A2(new_n767_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n247_), .B(new_n772_), .C1(new_n704_), .C2(new_n706_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n779_), .B(new_n783_), .C1(new_n784_), .C2(new_n513_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT112), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n783_), .C1(new_n784_), .C2(new_n513_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT51), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n684_), .B(new_n771_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n782_), .B1(new_n791_), .B2(G99gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n792_), .B2(new_n779_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n769_), .A2(new_n502_), .A3(new_n692_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n692_), .B(new_n771_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n796_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  NAND2_X1  g604(.A1(new_n486_), .A2(new_n622_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n597_), .A2(new_n598_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n808_), .A2(new_n591_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT12), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n599_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n809_), .A2(KEYINPUT55), .A3(new_n811_), .A4(new_n602_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n606_), .A2(KEYINPUT67), .A3(new_n607_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n610_), .B1(new_n609_), .B2(new_n522_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n600_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n524_), .A2(new_n526_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT12), .B1(new_n818_), .B2(new_n592_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n602_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n614_), .A2(new_n603_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n614_), .B2(new_n603_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n814_), .A2(new_n821_), .A3(new_n822_), .A4(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n619_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n619_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n807_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT117), .B(new_n807_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n469_), .A2(new_n470_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n462_), .A2(new_n470_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n485_), .B1(new_n833_), .B2(new_n479_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n481_), .A2(new_n485_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n623_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n831_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n660_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n665_), .A2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n825_), .A2(new_n619_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n619_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n806_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n836_), .B1(new_n846_), .B2(KEYINPUT117), .ZN(new_n847_));
  INV_X1    g646(.A(new_n831_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n841_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n844_), .A2(new_n845_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(KEYINPUT119), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n835_), .A2(new_n622_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n835_), .A2(new_n622_), .A3(KEYINPUT118), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n858_), .A2(new_n859_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n852_), .A2(new_n855_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n855_), .B1(new_n852_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n571_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n837_), .A2(KEYINPUT121), .A3(new_n841_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n840_), .A2(new_n851_), .A3(new_n865_), .A4(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n627_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n742_), .A2(new_n868_), .A3(new_n625_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n570_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT115), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n570_), .A2(new_n873_), .A3(new_n870_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n570_), .B2(new_n870_), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT115), .B(new_n869_), .C1(new_n562_), .C2(new_n569_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n867_), .A2(new_n643_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n667_), .A2(new_n438_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n419_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(G113gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n486_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n883_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n876_), .A2(new_n880_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n837_), .A2(KEYINPUT121), .A3(new_n841_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT121), .B1(new_n837_), .B2(new_n841_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n839_), .A2(new_n838_), .B1(new_n571_), .B2(new_n864_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n642_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT59), .B(new_n889_), .C1(new_n890_), .C2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n487_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n886_), .B1(new_n897_), .B2(new_n885_), .ZN(G1340gat));
  INV_X1    g697(.A(G120gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(KEYINPUT60), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n628_), .B2(KEYINPUT60), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(KEYINPUT122), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n884_), .B(new_n902_), .C1(KEYINPUT122), .C2(new_n901_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n628_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n899_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT123), .B(new_n903_), .C1(new_n904_), .C2(new_n899_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1341gat));
  INV_X1    g708(.A(G127gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n884_), .A2(new_n910_), .A3(new_n642_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n643_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(G1342gat));
  INV_X1    g712(.A(G134gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n884_), .A2(new_n914_), .A3(new_n665_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n570_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n914_), .ZN(G1343gat));
  NOR2_X1   g716(.A1(new_n881_), .A2(new_n433_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n882_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n487_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT124), .B(G141gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1344gat));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n629_), .A3(new_n882_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g723(.A1(new_n919_), .A2(new_n643_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT61), .B(G155gat), .Z(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n919_), .B2(new_n570_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n665_), .A2(new_n255_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n919_), .B2(new_n929_), .ZN(G1347gat));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n867_), .A2(new_n643_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n876_), .A2(new_n880_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n655_), .A2(new_n352_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n934_), .A2(new_n419_), .A3(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n487_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n931_), .B1(new_n937_), .B2(new_n205_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT62), .B(G169gat), .C1(new_n936_), .C2(new_n487_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n357_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(G1348gat));
  OR2_X1    g740(.A1(new_n936_), .A2(new_n628_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n206_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n225_), .B2(new_n942_), .ZN(G1349gat));
  NOR2_X1   g743(.A1(new_n936_), .A2(new_n643_), .ZN(new_n945_));
  MUX2_X1   g744(.A(G183gat), .B(new_n210_), .S(new_n945_), .Z(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n936_), .B2(new_n570_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n665_), .A2(new_n211_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n936_), .B2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(KEYINPUT125), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n947_), .B(new_n951_), .C1(new_n936_), .C2(new_n948_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(G1351gat));
  AND3_X1   g752(.A1(new_n934_), .A2(new_n434_), .A3(new_n935_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n486_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n629_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n642_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n959_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT63), .B(G211gat), .Z(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n959_), .B2(new_n961_), .ZN(G1354gat));
  NAND2_X1  g761(.A1(new_n918_), .A2(new_n935_), .ZN(new_n963_));
  OAI21_X1  g762(.A(G218gat), .B1(new_n963_), .B2(new_n570_), .ZN(new_n964_));
  INV_X1    g763(.A(G218gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n665_), .A2(new_n965_), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n964_), .B(KEYINPUT126), .C1(new_n963_), .C2(new_n966_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n965_), .B1(new_n954_), .B2(new_n571_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n963_), .A2(new_n966_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n968_), .B1(new_n969_), .B2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n967_), .A2(new_n971_), .ZN(G1355gat));
endmodule


