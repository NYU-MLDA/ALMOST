//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n203_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(G141gat), .C2(G148gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n204_), .B(new_n205_), .C1(KEYINPUT84), .C2(KEYINPUT3), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  AND3_X1   g014(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n213_), .A2(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n218_), .A2(KEYINPUT85), .B1(new_n207_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n202_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n210_), .B1(new_n223_), .B2(KEYINPUT86), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n202_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT28), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n224_), .A2(new_n231_), .A3(new_n225_), .A4(new_n228_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G22gat), .B(G50gat), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G78gat), .B(G106gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n223_), .A2(KEYINPUT86), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n203_), .A2(new_n209_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT29), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G228gat), .ZN(new_n243_));
  INV_X1    g042(.A(G233gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(G197gat), .A2(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(KEYINPUT21), .A3(new_n248_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n242_), .A2(new_n246_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n246_), .B1(new_n242_), .B2(new_n259_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n237_), .B(new_n238_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n225_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n257_), .A2(new_n258_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n245_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n242_), .A2(new_n246_), .A3(new_n259_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n238_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n266_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n237_), .B1(new_n270_), .B2(new_n238_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n236_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G113gat), .B(G120gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n273_), .A2(new_n274_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G43gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n281_), .A2(G43gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT30), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(G15gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n281_), .A2(G43gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n282_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n285_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n285_), .B2(new_n291_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT79), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G183gat), .A3(G190gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT23), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n301_));
  INV_X1    g100(.A(new_n296_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G183gat), .ZN(new_n306_));
  INV_X1    g105(.A(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n297_), .A2(new_n299_), .A3(new_n301_), .A4(KEYINPUT23), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT78), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(KEYINPUT24), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT25), .B(G183gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G190gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n320_), .A2(new_n321_), .B1(new_n322_), .B2(new_n317_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n302_), .A2(new_n303_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT23), .B1(new_n297_), .B2(new_n299_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n319_), .B(new_n323_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n316_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT82), .B1(new_n295_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n316_), .A2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n280_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT82), .ZN(new_n332_));
  INV_X1    g131(.A(new_n294_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n333_), .A3(new_n292_), .ZN(new_n334_));
  AND4_X1   g133(.A1(new_n332_), .A2(new_n334_), .A3(new_n280_), .A4(new_n330_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n279_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n332_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n330_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT31), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(new_n280_), .A3(new_n330_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n279_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n238_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT89), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n234_), .A2(new_n235_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n270_), .A2(new_n347_), .A3(new_n238_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .A4(new_n268_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n272_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n354_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n352_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n351_), .A3(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT97), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n364_), .A3(KEYINPUT97), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372_));
  INV_X1    g171(.A(G169gat), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n373_), .A2(KEYINPUT22), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(KEYINPUT22), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n372_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n311_), .A2(KEYINPUT90), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n312_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n308_), .B1(new_n325_), .B2(new_n324_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n315_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n318_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n323_), .A2(new_n305_), .A3(new_n309_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT20), .B1(new_n383_), .B2(new_n259_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n316_), .A2(new_n326_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n371_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n259_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n316_), .A2(new_n326_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n371_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(KEYINPUT20), .A4(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n369_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n388_), .A3(KEYINPUT20), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n371_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n329_), .A2(new_n259_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n264_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT20), .A4(new_n389_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n393_), .A2(new_n365_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n391_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n365_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT98), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT98), .B(new_n398_), .C1(new_n397_), .C2(new_n400_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G85gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT0), .B(G57gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n279_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n223_), .A2(KEYINPUT86), .ZN(new_n412_));
  INV_X1    g211(.A(new_n278_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n275_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(new_n228_), .A3(new_n240_), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(KEYINPUT4), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n279_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n416_), .A2(KEYINPUT93), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n420_), .A2(new_n418_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT93), .B1(new_n424_), .B2(new_n416_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n410_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT93), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n411_), .A2(KEYINPUT4), .A3(new_n415_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n418_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n430_), .A2(new_n409_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n426_), .A2(KEYINPUT96), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT96), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n433_), .B(new_n410_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n350_), .A2(new_n405_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n350_), .A2(new_n405_), .A3(KEYINPUT99), .A4(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n343_), .B(KEYINPUT83), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n272_), .A2(new_n349_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n405_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n443_));
  AND4_X1   g242(.A1(KEYINPUT32), .A2(new_n386_), .A3(new_n365_), .A4(new_n390_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n393_), .A2(new_n396_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(KEYINPUT95), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT95), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n432_), .A2(new_n450_), .A3(new_n434_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n423_), .A2(new_n425_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT94), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n409_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n431_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n365_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n445_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n416_), .A2(new_n417_), .A3(new_n420_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n411_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n410_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n393_), .A2(new_n365_), .A3(new_n396_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n459_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n442_), .B1(new_n451_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n441_), .B1(new_n443_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n440_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G29gat), .B(G36gat), .Z(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G8gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT74), .ZN(new_n476_));
  INV_X1    g275(.A(G22gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n287_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G15gat), .A2(G22gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G1gat), .A2(G8gat), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n478_), .A2(new_n479_), .B1(KEYINPUT14), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n476_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n471_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n474_), .B1(new_n484_), .B2(new_n473_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G229gat), .A2(G233gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n484_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT77), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n489_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n495_));
  OR2_X1    g294(.A1(G85gat), .A2(G92gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT7), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n501_), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n508_), .B(new_n507_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(KEYINPUT64), .A3(new_n498_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(KEYINPUT8), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n500_), .A2(new_n502_), .ZN(new_n518_));
  OR2_X1    g317(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n506_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n496_), .A2(KEYINPUT9), .A3(new_n497_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n497_), .A2(KEYINPUT9), .ZN(new_n523_));
  AND4_X1   g322(.A1(new_n518_), .A2(new_n521_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT64), .B1(new_n515_), .B2(new_n498_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(G78gat), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  INV_X1    g331(.A(G78gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n528_), .ZN(new_n534_));
  INV_X1    g333(.A(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G57gat), .ZN(new_n536_));
  INV_X1    g335(.A(G57gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G64gat), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n538_), .A3(KEYINPUT11), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT11), .B1(new_n536_), .B2(new_n538_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n531_), .B(new_n534_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n538_), .A3(KEYINPUT11), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n533_), .B1(new_n532_), .B2(new_n528_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n529_), .A2(new_n530_), .A3(G78gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n541_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n517_), .B(new_n527_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT68), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n547_), .A2(new_n548_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n517_), .A2(new_n527_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT12), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n517_), .A2(new_n527_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n517_), .B2(new_n527_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n558_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n555_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n556_), .A2(new_n557_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n549_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(G230gat), .A3(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n566_), .A2(new_n569_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n573_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n575_), .A2(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT70), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n586_), .B2(new_n578_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n495_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n582_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n584_), .A3(new_n578_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(KEYINPUT13), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n494_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n468_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n517_), .A2(new_n527_), .A3(new_n559_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n471_), .B(new_n472_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n517_), .A2(new_n527_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n471_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n597_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n604_), .A3(new_n597_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT72), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n601_), .A2(new_n604_), .A3(new_n597_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n605_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(new_n610_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n615_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n610_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT73), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n594_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n621_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT37), .B(new_n626_), .C1(new_n613_), .C2(new_n617_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n482_), .B(new_n629_), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n541_), .A2(new_n545_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT75), .Z(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634_));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635_));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n633_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n630_), .B(new_n556_), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n639_), .B(KEYINPUT17), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n628_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n593_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT100), .Z(new_n648_));
  INV_X1    g447(.A(G1gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n435_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n648_), .A2(KEYINPUT38), .A3(new_n649_), .A4(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n468_), .A2(new_n592_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n626_), .B1(new_n613_), .B2(new_n617_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n655_), .A2(new_n645_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n435_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n654_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n653_), .A2(KEYINPUT101), .A3(new_n654_), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(G8gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n405_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n657_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT39), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n648_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(new_n441_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n287_), .B1(new_n657_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n287_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n647_), .B2(new_n676_), .ZN(G1326gat));
  AOI21_X1  g476(.A(new_n477_), .B1(new_n657_), .B2(new_n442_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT42), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n442_), .A2(new_n477_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT102), .Z(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n647_), .B2(new_n681_), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n656_), .A2(new_n645_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT105), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n468_), .A2(new_n592_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT106), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n468_), .A2(new_n592_), .A3(new_n684_), .A4(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n650_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n592_), .A2(new_n645_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n405_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n451_), .A2(new_n465_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n442_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n694_), .A2(new_n441_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n656_), .A2(new_n594_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n613_), .A2(new_n617_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n696_), .B(new_n697_), .C1(new_n698_), .C2(new_n594_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n624_), .B2(new_n627_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n695_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n628_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n440_), .B2(new_n467_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n691_), .B1(new_n702_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT44), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n589_), .A2(new_n590_), .A3(KEYINPUT13), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT13), .B1(new_n589_), .B2(new_n590_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n645_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n711_), .A2(new_n494_), .A3(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n699_), .A2(new_n700_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n703_), .B1(new_n468_), .B2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT44), .B(new_n713_), .C1(new_n715_), .C2(new_n705_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n717_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n708_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n650_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n690_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n405_), .A2(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n686_), .A2(new_n688_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT107), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n686_), .A2(new_n728_), .A3(new_n688_), .A4(new_n725_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n727_), .A2(KEYINPUT45), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n727_), .B2(new_n729_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n702_), .A2(new_n706_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n713_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT104), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n666_), .B(new_n736_), .C1(new_n737_), .C2(new_n718_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G36gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n724_), .B1(new_n732_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n732_), .A2(new_n739_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT109), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1329gat));
  AOI21_X1  g544(.A(G43gat), .B1(new_n689_), .B2(new_n673_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n343_), .A2(G43gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n721_), .B2(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g548(.A(G50gat), .B1(new_n689_), .B2(new_n442_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n442_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n721_), .B2(new_n751_), .ZN(G1331gat));
  NAND2_X1  g551(.A1(new_n588_), .A2(new_n591_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n494_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n468_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n756_), .A2(new_n645_), .A3(new_n656_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n435_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n756_), .A2(new_n645_), .A3(new_n628_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n537_), .A3(new_n650_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1332gat));
  AOI21_X1  g561(.A(new_n535_), .B1(new_n757_), .B2(new_n666_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT48), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n535_), .A3(new_n666_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n757_), .B2(new_n673_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n767_), .A3(new_n673_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1334gat));
  AOI21_X1  g570(.A(new_n533_), .B1(new_n757_), .B2(new_n442_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n760_), .A2(new_n533_), .A3(new_n442_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1335gat));
  OR2_X1    g575(.A1(new_n733_), .A2(KEYINPUT111), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n733_), .A2(KEYINPUT111), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n753_), .A2(new_n754_), .A3(new_n712_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT112), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n777_), .A2(new_n778_), .A3(new_n782_), .A4(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n435_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n755_), .A2(new_n468_), .A3(new_n684_), .ZN(new_n786_));
  INV_X1    g585(.A(G85gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n650_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n786_), .B2(new_n666_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT113), .Z(new_n791_));
  NAND2_X1  g590(.A1(new_n666_), .A2(G92gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n784_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT114), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n791_), .C1(new_n784_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1337gat));
  NAND4_X1  g596(.A1(new_n786_), .A2(new_n519_), .A3(new_n520_), .A4(new_n343_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n777_), .A2(new_n778_), .A3(new_n673_), .A4(new_n779_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n799_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT115), .B1(new_n799_), .B2(G99gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT51), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n798_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1338gat));
  AND3_X1   g605(.A1(new_n733_), .A2(new_n442_), .A3(new_n779_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n807_), .A2(KEYINPUT52), .A3(new_n506_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n807_), .B2(new_n506_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n786_), .A2(new_n506_), .A3(new_n442_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1339gat));
  NAND2_X1  g613(.A1(new_n350_), .A2(new_n405_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n493_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n485_), .A2(new_n486_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n488_), .B2(new_n486_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n489_), .A2(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n575_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n598_), .A2(new_n599_), .A3(new_n564_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n567_), .A2(new_n563_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n549_), .ZN(new_n825_));
  OAI211_X1 g624(.A(G230gat), .B(G233gat), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n555_), .B2(new_n565_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n826_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n549_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n553_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT117), .B1(new_n833_), .B2(new_n824_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(KEYINPUT55), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n573_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(KEYINPUT55), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n828_), .A2(new_n829_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n826_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT56), .A3(new_n573_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n821_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n628_), .B1(new_n843_), .B2(KEYINPUT58), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n845_), .B(new_n821_), .C1(new_n838_), .C2(new_n842_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n656_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n754_), .A2(new_n575_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n550_), .B1(new_n565_), .B2(new_n549_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n834_), .B2(KEYINPUT55), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n837_), .B(new_n574_), .C1(new_n851_), .C2(new_n840_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n838_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n841_), .B2(new_n573_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT118), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n849_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n589_), .A2(new_n590_), .A3(new_n820_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n848_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n847_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n754_), .A2(new_n575_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n842_), .B1(new_n855_), .B2(KEYINPUT118), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n838_), .A2(new_n853_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n858_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n656_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT57), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n712_), .B1(new_n861_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n696_), .B1(new_n594_), .B2(new_n698_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n494_), .A3(new_n712_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n711_), .A2(KEYINPUT54), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873_));
  INV_X1    g672(.A(new_n871_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n753_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n650_), .B(new_n816_), .C1(new_n869_), .C2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(G113gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n754_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n881_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n844_), .A2(new_n846_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n867_), .B2(KEYINPUT57), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n859_), .A2(new_n860_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n645_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n876_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(KEYINPUT59), .A3(new_n650_), .A4(new_n816_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n494_), .B1(new_n882_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n880_), .B1(new_n890_), .B2(new_n879_), .ZN(G1340gat));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n753_), .B2(KEYINPUT60), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(KEYINPUT60), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(KEYINPUT119), .B2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n878_), .B(new_n895_), .C1(KEYINPUT119), .C2(new_n893_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n753_), .B1(new_n882_), .B2(new_n889_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  OAI21_X1  g697(.A(G120gat), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n435_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT59), .B1(new_n900_), .B2(new_n816_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n838_), .A2(new_n853_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n856_), .A3(new_n842_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n858_), .B1(new_n903_), .B2(new_n862_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n860_), .B1(new_n904_), .B2(new_n656_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n868_), .A2(new_n905_), .A3(new_n883_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n876_), .B1(new_n906_), .B2(new_n645_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n907_), .A2(new_n881_), .A3(new_n435_), .A4(new_n815_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n898_), .B(new_n711_), .C1(new_n901_), .C2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n896_), .B1(new_n899_), .B2(new_n910_), .ZN(G1341gat));
  INV_X1    g710(.A(G127gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n878_), .A2(new_n912_), .A3(new_n712_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n645_), .B1(new_n882_), .B2(new_n889_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n912_), .ZN(G1342gat));
  INV_X1    g714(.A(G134gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n878_), .A2(new_n916_), .A3(new_n656_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n870_), .B1(new_n882_), .B2(new_n889_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1343gat));
  NAND3_X1  g718(.A1(new_n441_), .A2(new_n442_), .A3(new_n405_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n907_), .A2(new_n435_), .A3(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n754_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n711_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT121), .B(G148gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1345gat));
  NAND2_X1  g725(.A1(new_n921_), .A2(new_n712_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT122), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n921_), .A2(new_n929_), .A3(new_n712_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n928_), .A2(new_n930_), .A3(new_n932_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1346gat));
  NAND3_X1  g735(.A1(new_n921_), .A2(G162gat), .A3(new_n714_), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n907_), .A2(new_n435_), .A3(new_n848_), .A4(new_n920_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(G162gat), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n937_), .B(KEYINPUT123), .C1(new_n938_), .C2(G162gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1347gat));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n441_), .A2(new_n650_), .A3(new_n405_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  NOR4_X1   g745(.A1(new_n907_), .A2(new_n494_), .A3(new_n442_), .A4(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  OAI21_X1  g749(.A(G169gat), .B1(new_n947_), .B2(new_n948_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n944_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n907_), .A2(new_n442_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n945_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT124), .B1(new_n954_), .B2(new_n494_), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n955_), .A2(KEYINPUT62), .A3(new_n949_), .A4(G169gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n947_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n952_), .A2(new_n956_), .A3(new_n957_), .ZN(G1348gat));
  INV_X1    g757(.A(new_n954_), .ZN(new_n959_));
  AOI21_X1  g758(.A(G176gat), .B1(new_n959_), .B2(new_n711_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n953_), .B(KEYINPUT125), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n753_), .A2(new_n946_), .A3(new_n312_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n960_), .B1(new_n961_), .B2(new_n962_), .ZN(G1349gat));
  NOR3_X1   g762(.A1(new_n954_), .A2(new_n320_), .A3(new_n645_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n961_), .A2(new_n712_), .A3(new_n945_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n965_), .B2(new_n306_), .ZN(G1350gat));
  OAI21_X1  g765(.A(G190gat), .B1(new_n954_), .B2(new_n870_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n656_), .A2(new_n321_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n954_), .B2(new_n968_), .ZN(G1351gat));
  AND4_X1   g768(.A1(new_n441_), .A2(new_n442_), .A3(new_n435_), .A4(new_n666_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n888_), .A2(new_n970_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(new_n754_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g773(.A1(new_n971_), .A2(new_n753_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(G204gat), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n977_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(KEYINPUT126), .B(G204gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n975_), .B2(new_n979_), .ZN(G1353gat));
  AOI21_X1  g779(.A(new_n645_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n981_));
  INV_X1    g780(.A(new_n981_), .ZN(new_n982_));
  OR3_X1    g781(.A1(new_n971_), .A2(KEYINPUT127), .A3(new_n982_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n984_));
  OAI21_X1  g783(.A(KEYINPUT127), .B1(new_n971_), .B2(new_n982_), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n983_), .A2(new_n984_), .A3(new_n985_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n984_), .B1(new_n983_), .B2(new_n985_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1354gat));
  OR3_X1    g787(.A1(new_n971_), .A2(G218gat), .A3(new_n848_), .ZN(new_n989_));
  OAI21_X1  g788(.A(G218gat), .B1(new_n971_), .B2(new_n870_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n989_), .A2(new_n990_), .ZN(G1355gat));
endmodule


