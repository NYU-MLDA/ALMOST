//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n207_), .B(new_n208_), .Z(new_n209_));
  XOR2_X1   g008(.A(G29gat), .B(G36gat), .Z(new_n210_));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT76), .B1(new_n209_), .B2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n209_), .A2(new_n212_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G229gat), .A3(G233gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n212_), .B(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n218_), .A2(new_n209_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n209_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n212_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n219_), .B(new_n220_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G113gat), .B(G141gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G169gat), .B(G197gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n224_), .B(new_n225_), .Z(new_n226_));
  NAND3_X1  g025(.A1(new_n216_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n216_), .B2(new_n223_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n202_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT77), .A3(new_n227_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n239_));
  INV_X1    g038(.A(G169gat), .ZN(new_n240_));
  INV_X1    g039(.A(G176gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT24), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n244_), .ZN(new_n249_));
  INV_X1    g048(.A(G190gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT26), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT79), .ZN(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT25), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(KEYINPUT79), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n257_), .A2(G183gat), .B1(new_n258_), .B2(G190gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n252_), .A2(new_n255_), .A3(new_n256_), .A4(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G183gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT23), .B1(new_n261_), .B2(new_n250_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(G183gat), .A3(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n249_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n262_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n253_), .A2(new_n254_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n268_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n266_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n266_), .A2(KEYINPUT82), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281_));
  INV_X1    g080(.A(G43gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n280_), .B(new_n283_), .Z(new_n284_));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(G15gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT30), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n280_), .B(new_n283_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n238_), .B1(new_n292_), .B2(KEYINPUT84), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT84), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n288_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300_));
  INV_X1    g099(.A(G155gat), .ZN(new_n301_));
  INV_X1    g100(.A(G162gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT88), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n303_), .A2(new_n308_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT2), .Z(new_n311_));
  NOR2_X1   g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n307_), .B(new_n309_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n318_), .A2(new_n319_), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n305_), .A2(KEYINPUT1), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(G155gat), .A3(G162gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n303_), .A2(new_n321_), .A3(new_n323_), .A4(new_n304_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n315_), .B(new_n316_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n236_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n328_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n326_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n236_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n316_), .A3(new_n333_), .A4(new_n315_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n299_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT99), .B(KEYINPUT4), .Z(new_n336_));
  AOI211_X1 g135(.A(new_n236_), .B(new_n336_), .C1(new_n332_), .C2(new_n315_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n298_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  AND2_X1   g142(.A1(new_n330_), .A2(new_n334_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n297_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n338_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n343_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n292_), .A2(KEYINPUT84), .A3(new_n238_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n296_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352_));
  XOR2_X1   g151(.A(G8gat), .B(G36gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT19), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT94), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT92), .ZN(new_n363_));
  INV_X1    g162(.A(G204gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G197gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n368_));
  INV_X1    g167(.A(G197gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G204gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n361_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n363_), .A2(KEYINPUT21), .A3(new_n371_), .A4(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n367_), .A2(new_n368_), .A3(new_n375_), .A4(new_n370_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT91), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n362_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n376_), .A2(new_n377_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n374_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n278_), .A2(new_n384_), .A3(new_n279_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT25), .B(G183gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n258_), .A2(G190gat), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n387_), .A2(new_n251_), .A3(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n272_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n249_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n265_), .B1(G183gat), .B2(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n245_), .A2(KEYINPUT95), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n245_), .A2(KEYINPUT95), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G169gat), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n393_), .A2(new_n394_), .B1(new_n395_), .B2(new_n241_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n386_), .B1(new_n398_), .B2(new_n383_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n360_), .B1(new_n385_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n398_), .B2(new_n383_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n280_), .B2(new_n383_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n400_), .A2(new_n401_), .B1(new_n403_), .B2(new_n359_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n385_), .A2(new_n399_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n360_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT96), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n357_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n266_), .A2(KEYINPUT82), .A3(new_n275_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT82), .B1(new_n266_), .B2(new_n275_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n383_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n390_), .A2(new_n249_), .B1(new_n396_), .B2(new_n392_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n401_), .B(new_n406_), .C1(new_n412_), .C2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n383_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n386_), .B1(new_n384_), .B2(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n359_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n357_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n401_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n352_), .B1(new_n409_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT102), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n412_), .A2(new_n414_), .A3(new_n406_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n359_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n420_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT27), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n332_), .A2(new_n315_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT29), .ZN(new_n431_));
  AND2_X1   g230(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(G233gat), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n434_), .A3(new_n383_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n436_));
  AOI21_X1  g235(.A(new_n384_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n437_), .B2(new_n434_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G78gat), .B(G106gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT28), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n332_), .A2(new_n442_), .A3(new_n443_), .A4(new_n315_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G22gat), .B(G50gat), .Z(new_n445_));
  AND3_X1   g244(.A1(new_n441_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n439_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n435_), .B(new_n449_), .C1(new_n437_), .C2(new_n434_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n440_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n440_), .B2(new_n450_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n404_), .A2(new_n357_), .A3(new_n408_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n403_), .A2(new_n359_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n352_), .B1(new_n455_), .B2(new_n420_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n456_), .A3(KEYINPUT102), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n423_), .A2(new_n429_), .A3(new_n453_), .A4(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT103), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n351_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n420_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n454_), .A2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n347_), .A2(KEYINPUT33), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n335_), .A2(new_n298_), .A3(new_n337_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n343_), .B1(new_n344_), .B2(new_n297_), .ZN(new_n467_));
  OAI22_X1  g266(.A1(new_n347_), .A2(KEYINPUT33), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n464_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n425_), .A2(new_n426_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n357_), .A2(KEYINPUT32), .ZN(new_n471_));
  OAI22_X1  g270(.A1(new_n346_), .A2(new_n347_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n404_), .A2(new_n471_), .A3(new_n408_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT101), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT101), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n404_), .A2(new_n408_), .A3(new_n475_), .A4(new_n471_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n453_), .B1(new_n469_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n348_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n480_), .A2(new_n429_), .A3(new_n423_), .A4(new_n457_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n296_), .A2(new_n349_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n233_), .B1(new_n462_), .B2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(KEYINPUT66), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(KEYINPUT66), .A2(G106gat), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(G85gat), .A2(G92gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT9), .ZN(new_n493_));
  AND2_X1   g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT67), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n492_), .B(new_n493_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT6), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n492_), .A2(KEYINPUT67), .A3(KEYINPUT9), .A4(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n491_), .A2(new_n496_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  INV_X1    g305(.A(new_n490_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n486_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n506_), .A2(new_n508_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n496_), .A4(new_n503_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  OR3_X1    g311(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n501_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n494_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT8), .B1(new_n516_), .B2(KEYINPUT69), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n514_), .A2(new_n517_), .A3(new_n516_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n516_), .B2(new_n514_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n505_), .B(new_n511_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n521_));
  INV_X1    g320(.A(G71gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G78gat), .ZN(new_n523_));
  INV_X1    g322(.A(G78gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G71gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(KEYINPUT11), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n527_), .B2(KEYINPUT11), .ZN(new_n530_));
  INV_X1    g329(.A(G64gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(G57gat), .ZN(new_n532_));
  INV_X1    g331(.A(G57gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(G64gat), .ZN(new_n534_));
  AND4_X1   g333(.A1(new_n529_), .A2(new_n532_), .A3(new_n534_), .A4(KEYINPUT11), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n528_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n534_), .A3(KEYINPUT11), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT70), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n534_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT11), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n532_), .A2(new_n534_), .A3(new_n529_), .A4(KEYINPUT11), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n538_), .A2(new_n541_), .A3(new_n526_), .A4(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n521_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n520_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(new_n543_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n536_), .A2(new_n543_), .A3(KEYINPUT71), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n545_), .B1(new_n550_), .B2(new_n520_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT12), .B1(new_n550_), .B2(new_n520_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n551_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n520_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n518_), .A2(new_n519_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n511_), .A2(new_n505_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n548_), .A4(new_n549_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NOR3_X1   g365(.A1(new_n556_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n218_), .A2(new_n520_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n559_), .A2(new_n560_), .A3(new_n222_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n581_), .B1(KEYINPUT73), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  XOR2_X1   g387(.A(G134gat), .B(G162gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n586_), .A2(KEYINPUT73), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n587_), .A2(new_n588_), .A3(new_n591_), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n588_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n591_), .A2(new_n588_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n577_), .A2(new_n584_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n597_), .A2(new_n598_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n595_), .B(new_n596_), .C1(new_n599_), .C2(new_n592_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(new_n603_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT17), .Z(new_n611_));
  INV_X1    g410(.A(new_n550_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n209_), .B(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n614_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n614_), .A2(new_n546_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n546_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n618_), .A2(KEYINPUT17), .A3(new_n619_), .A4(new_n610_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n604_), .A2(new_n605_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n485_), .A2(new_n574_), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT104), .ZN(new_n624_));
  INV_X1    g423(.A(new_n348_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n204_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n594_), .A2(new_n600_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT105), .Z(new_n630_));
  AOI211_X1 g429(.A(new_n621_), .B(new_n630_), .C1(new_n462_), .C2(new_n484_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n574_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(new_n233_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n348_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n626_), .A2(new_n627_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  AND3_X1   g436(.A1(new_n454_), .A2(new_n456_), .A3(KEYINPUT102), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT27), .B1(new_n454_), .B2(new_n463_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n429_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n624_), .A2(new_n205_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n631_), .A2(new_n641_), .A3(new_n633_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(G8gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n643_), .A3(G8gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n634_), .B2(new_n483_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT41), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n623_), .A2(G15gat), .A3(new_n483_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  OAI21_X1  g453(.A(G22gat), .B1(new_n634_), .B2(new_n453_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT42), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n453_), .A2(G22gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n623_), .B2(new_n657_), .ZN(G1327gat));
  NAND3_X1  g457(.A1(new_n594_), .A2(new_n600_), .A3(new_n621_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n632_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n485_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n625_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n462_), .A2(new_n484_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n602_), .B(KEYINPUT37), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .A4(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n640_), .A2(KEYINPUT103), .A3(new_n453_), .A4(new_n429_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n458_), .A2(new_n459_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n350_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n292_), .A2(KEYINPUT84), .A3(new_n238_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n666_), .B(new_n668_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT107), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n668_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT43), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n669_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n621_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n632_), .A2(new_n233_), .A3(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT106), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT44), .B1(new_n680_), .B2(new_n683_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n625_), .A2(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n663_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(new_n641_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n661_), .A2(G36gat), .A3(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT45), .Z(new_n691_));
  NOR3_X1   g490(.A1(new_n684_), .A2(new_n685_), .A3(new_n689_), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT46), .B(new_n691_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1329gat));
  NOR2_X1   g497(.A1(new_n483_), .A2(new_n282_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n686_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G43gat), .B1(new_n662_), .B2(new_n674_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n700_), .A2(new_n702_), .A3(new_n704_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1330gat));
  INV_X1    g507(.A(new_n453_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G50gat), .B1(new_n662_), .B2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n686_), .B2(new_n711_), .ZN(G1331gat));
  INV_X1    g511(.A(new_n233_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n574_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n631_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n348_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n462_), .B2(new_n484_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n622_), .A2(new_n632_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n533_), .A3(new_n625_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n715_), .B2(new_n689_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n641_), .A2(new_n531_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT109), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n719_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n715_), .B2(new_n483_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n720_), .A2(new_n522_), .A3(new_n674_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1334gat));
  NAND3_X1  g530(.A1(new_n720_), .A2(new_n524_), .A3(new_n709_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n631_), .A2(new_n709_), .A3(new_n714_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(G78gat), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n733_), .B2(G78gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT111), .Z(G1335gat));
  NOR3_X1   g538(.A1(new_n574_), .A2(new_n713_), .A3(new_n681_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n680_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n348_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n574_), .A2(new_n659_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n717_), .A2(new_n743_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n744_), .A2(G85gat), .A3(new_n348_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1336gat));
  INV_X1    g545(.A(new_n744_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G92gat), .B1(new_n747_), .B2(new_n641_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n741_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n641_), .A2(G92gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT112), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n749_), .B2(new_n751_), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n741_), .B2(new_n483_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n674_), .A3(new_n506_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n754_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n709_), .A3(new_n508_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n680_), .A2(new_n709_), .A3(new_n740_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n762_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  XNOR2_X1  g570(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n667_), .A2(new_n574_), .A3(new_n681_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n713_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n622_), .A2(new_n233_), .A3(new_n574_), .A4(new_n772_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n215_), .A2(new_n220_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n220_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n226_), .B1(new_n219_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n227_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n567_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n559_), .A2(new_n560_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n561_), .B(new_n545_), .C1(new_n787_), .C2(KEYINPUT12), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n785_), .B(new_n786_), .C1(new_n788_), .C2(new_n555_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n788_), .B2(new_n555_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n790_), .B(new_n555_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n556_), .A2(KEYINPUT55), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n551_), .A2(new_n552_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(new_n796_), .B2(new_n557_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n785_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n566_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n555_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n792_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n556_), .B2(KEYINPUT55), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n795_), .A4(new_n789_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n784_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT58), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n566_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n783_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(KEYINPUT118), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n668_), .A3(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n230_), .A2(new_n232_), .A3(new_n568_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n570_), .A2(new_n782_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n629_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT57), .B(new_n629_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n777_), .B1(new_n621_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n348_), .B(new_n483_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n816_), .A2(new_n822_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n816_), .A2(new_n822_), .A3(KEYINPUT119), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n823_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n777_), .B1(new_n834_), .B2(new_n621_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n827_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n829_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n233_), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n828_), .A2(G113gat), .A3(new_n233_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n838_), .B2(new_n574_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n574_), .A2(KEYINPUT60), .ZN(new_n843_));
  MUX2_X1   g642(.A(new_n843_), .B(KEYINPUT60), .S(G120gat), .Z(new_n844_));
  NAND3_X1  g643(.A1(new_n826_), .A2(new_n827_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n845_), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n838_), .B2(new_n621_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n828_), .A2(G127gat), .A3(new_n621_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1342gat));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n667_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n829_), .B(new_n851_), .C1(new_n835_), .C2(new_n837_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n630_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n850_), .B1(new_n828_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT120), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n850_), .C1(new_n828_), .C2(new_n853_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n852_), .A2(new_n855_), .A3(new_n857_), .ZN(G1343gat));
  NOR3_X1   g657(.A1(new_n674_), .A2(new_n453_), .A3(new_n348_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n826_), .A2(new_n689_), .A3(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n233_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n574_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g663(.A1(new_n860_), .A2(new_n621_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  OAI21_X1  g666(.A(G162gat), .B1(new_n860_), .B2(new_n667_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n630_), .A2(new_n302_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n860_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n689_), .A2(new_n350_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n823_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n681_), .B1(new_n873_), .B2(new_n833_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n453_), .B(new_n871_), .C1(new_n874_), .C2(new_n777_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n713_), .A3(new_n395_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n871_), .A2(new_n713_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n453_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n813_), .A2(KEYINPUT118), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n667_), .B1(new_n883_), .B2(KEYINPUT58), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n884_), .A2(new_n815_), .B1(new_n821_), .B2(new_n820_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n823_), .B1(new_n885_), .B2(KEYINPUT119), .ZN(new_n886_));
  INV_X1    g685(.A(new_n833_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n621_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n777_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n882_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n240_), .B1(new_n890_), .B2(KEYINPUT122), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n835_), .B2(new_n882_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n878_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n882_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n895_), .B(KEYINPUT122), .C1(new_n874_), .C2(new_n777_), .ZN(new_n896_));
  AND4_X1   g695(.A1(new_n878_), .A2(new_n893_), .A3(G169gat), .A4(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n877_), .B1(new_n894_), .B2(new_n897_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n876_), .B2(new_n632_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n871_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n681_), .B1(new_n885_), .B2(new_n823_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n453_), .B1(new_n901_), .B2(new_n777_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT123), .B(new_n453_), .C1(new_n901_), .C2(new_n777_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n574_), .A2(new_n241_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n899_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  OAI21_X1  g707(.A(new_n903_), .B1(new_n825_), .B2(new_n709_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n909_), .A2(new_n905_), .A3(new_n681_), .A4(new_n871_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT124), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n904_), .A2(new_n912_), .A3(new_n681_), .A4(new_n905_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n273_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n875_), .A2(new_n387_), .A3(new_n621_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n875_), .B2(new_n667_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n630_), .A2(new_n251_), .A3(new_n388_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n875_), .B2(new_n918_), .ZN(G1351gat));
  NOR3_X1   g718(.A1(new_n689_), .A2(new_n479_), .A3(new_n674_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n826_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n233_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n369_), .ZN(G1352gat));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n574_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n364_), .ZN(G1353gat));
  INV_X1    g724(.A(new_n921_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT125), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT126), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n928_), .B(new_n931_), .ZN(G1354gat));
  AND3_X1   g731(.A1(new_n926_), .A2(G218gat), .A3(new_n668_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n921_), .A2(new_n853_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n934_), .A2(KEYINPUT127), .ZN(new_n935_));
  AOI21_X1  g734(.A(G218gat), .B1(new_n934_), .B2(KEYINPUT127), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(G1355gat));
endmodule


