//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT82), .Z(new_n210_));
  OR2_X1    g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n210_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT84), .B(G176gat), .Z(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  OAI21_X1  g016(.A(G169gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(G169gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n218_), .C1(new_n216_), .C2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n225_), .B(new_n213_), .C1(new_n210_), .C2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT30), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT87), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n208_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n231_), .B2(new_n208_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G120gat), .Z(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT31), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT88), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G197gat), .B(G204gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT21), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G197gat), .B(G204gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT21), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n248_), .A2(new_n251_), .A3(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT3), .Z(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT2), .Z(new_n264_));
  OAI211_X1 g063(.A(new_n258_), .B(new_n260_), .C1(new_n262_), .C2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(KEYINPUT1), .B2(new_n258_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(KEYINPUT1), .B2(new_n258_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n261_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n263_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n257_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n245_), .B1(new_n256_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT90), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(KEYINPUT90), .B(new_n245_), .C1(new_n256_), .C2(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n254_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n270_), .A2(new_n245_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n282_), .A3(new_n278_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n265_), .A2(new_n269_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n257_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G22gat), .B(G50gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT28), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n289_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n284_), .B1(new_n286_), .B2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n281_), .A2(new_n285_), .A3(new_n283_), .A4(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT19), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT92), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n215_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n214_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n209_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n225_), .B(new_n213_), .C1(new_n303_), .C2(new_n226_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n256_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT20), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n228_), .B2(new_n254_), .ZN(new_n309_));
  AOI211_X1 g108(.A(KEYINPUT98), .B(new_n298_), .C1(new_n307_), .C2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n254_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n254_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT93), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT93), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n305_), .A2(new_n314_), .A3(new_n254_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n311_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n298_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT98), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n307_), .A2(new_n309_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n297_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n310_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G8gat), .B(G36gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n287_), .A2(new_n237_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n287_), .A2(new_n237_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(KEYINPUT4), .A3(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(KEYINPUT4), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G1gat), .B(G29gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n336_), .A2(new_n344_), .A3(new_n338_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n321_), .A2(new_n328_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n313_), .A2(new_n315_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n311_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT94), .A3(new_n297_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n316_), .B2(new_n298_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n306_), .A2(new_n276_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n309_), .A3(new_n298_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n357_), .A3(new_n327_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n294_), .A2(new_n295_), .B1(new_n348_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n326_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n326_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n357_), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n361_), .B(new_n362_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n346_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n331_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n329_), .A2(new_n335_), .A3(new_n330_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n344_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT97), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n367_), .A2(new_n368_), .A3(KEYINPUT97), .A4(new_n344_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n339_), .A2(KEYINPUT33), .A3(new_n345_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n366_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n242_), .B1(new_n359_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n346_), .A2(new_n347_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n321_), .B2(new_n361_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n355_), .A2(new_n326_), .A3(new_n357_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n294_), .A2(new_n295_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n377_), .A2(new_n387_), .A3(KEYINPUT99), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT99), .B1(new_n377_), .B2(new_n387_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n379_), .A2(new_n383_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n385_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n242_), .A2(new_n380_), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n388_), .A2(new_n389_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G57gat), .B(G64gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT11), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT67), .ZN(new_n396_));
  XOR2_X1   g195(.A(G71gat), .B(G78gat), .Z(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(KEYINPUT11), .B2(new_n394_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n396_), .B(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n400_));
  INV_X1    g199(.A(G106gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT64), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT64), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n400_), .A2(new_n405_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT66), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(G99gat), .B2(G106gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G99gat), .A2(G106gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(KEYINPUT6), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(KEYINPUT6), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(G99gat), .A3(G106gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT66), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G85gat), .A2(G92gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G85gat), .A2(G92gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n420_), .B2(KEYINPUT9), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT9), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT65), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n419_), .A2(KEYINPUT65), .A3(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n407_), .A2(new_n417_), .A3(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n420_), .A2(new_n418_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT8), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n429_), .B1(new_n417_), .B2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n432_), .B(new_n433_), .C1(new_n410_), .C2(new_n412_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n428_), .B1(new_n436_), .B2(new_n427_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n426_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n399_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n399_), .A2(new_n438_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G230gat), .A2(G233gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT66), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT66), .B1(new_n414_), .B2(new_n415_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n434_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n428_), .A3(new_n427_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n436_), .A2(new_n427_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT8), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(KEYINPUT68), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n445_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n426_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(KEYINPUT12), .A3(new_n399_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n442_), .A2(new_n443_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n439_), .ZN(new_n457_));
  OAI211_X1 g256(.A(G230gat), .B(G233gat), .C1(new_n457_), .C2(new_n440_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G120gat), .B(G148gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT5), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G176gat), .B(G204gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n459_), .A2(new_n464_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT13), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT78), .B(G15gat), .ZN(new_n473_));
  INV_X1    g272(.A(G22gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT79), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n481_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G36gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G29gat), .ZN(new_n486_));
  INV_X1    g285(.A(G29gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G36gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n486_), .A2(new_n488_), .A3(KEYINPUT70), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT70), .B1(new_n486_), .B2(new_n488_), .ZN(new_n490_));
  INV_X1    g289(.A(G50gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G43gat), .ZN(new_n492_));
  INV_X1    g291(.A(G43gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G50gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n489_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n492_), .A2(new_n494_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT70), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n487_), .A2(G36gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n485_), .A2(G29gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n486_), .A2(new_n488_), .A3(KEYINPUT70), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n497_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n484_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n495_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n502_), .A3(new_n497_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n508_), .A2(KEYINPUT15), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT15), .B1(new_n508_), .B2(new_n509_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n484_), .A2(new_n504_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n507_), .B(KEYINPUT81), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI22_X1  g317(.A1(new_n506_), .A2(new_n507_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G113gat), .B(G141gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G169gat), .B(G197gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n523_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n472_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n393_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n454_), .A2(KEYINPUT71), .A3(new_n513_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n531_));
  INV_X1    g330(.A(new_n426_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n533_), .B2(new_n512_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n504_), .B(new_n426_), .C1(new_n435_), .C2(new_n437_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n539_), .A2(new_n540_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n535_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n536_), .A2(KEYINPUT72), .A3(new_n541_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n534_), .B2(new_n530_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n543_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n551_), .A2(KEYINPUT73), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n554_));
  INV_X1    g353(.A(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT72), .B1(new_n536_), .B2(new_n541_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT71), .B1(new_n454_), .B2(new_n513_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n533_), .A2(new_n531_), .A3(new_n512_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n554_), .B1(new_n560_), .B2(new_n543_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n546_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G190gat), .B(G218gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT74), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT75), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n562_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT37), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n566_), .B(KEYINPUT36), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n562_), .A2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT73), .B1(new_n551_), .B2(new_n552_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n560_), .A2(new_n554_), .A3(new_n543_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n576_), .B1(new_n579_), .B2(new_n546_), .ZN(new_n580_));
  AOI211_X1 g379(.A(KEYINPUT76), .B(new_n545_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n573_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT77), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT77), .B(new_n573_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n570_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n575_), .B1(new_n586_), .B2(KEYINPUT37), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n484_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n399_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n597_), .B2(KEYINPUT17), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(KEYINPUT80), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT80), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n599_), .A3(new_n598_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n587_), .A2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n529_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n380_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n476_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n584_), .A2(new_n585_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT101), .B1(new_n613_), .B2(new_n571_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n615_), .B(new_n570_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n393_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n528_), .A2(new_n605_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT100), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n380_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n610_), .A2(new_n611_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n612_), .A2(new_n622_), .A3(new_n623_), .ZN(G1324gat));
  OAI21_X1  g423(.A(G8gat), .B1(new_n621_), .B2(new_n390_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT102), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n628_), .B(G8gat), .C1(new_n621_), .C2(new_n390_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(KEYINPUT39), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n390_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n608_), .A2(new_n477_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n627_), .A2(KEYINPUT40), .A3(new_n630_), .A4(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(new_n242_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G15gat), .B1(new_n621_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT41), .Z(new_n640_));
  INV_X1    g439(.A(G15gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n608_), .A2(new_n641_), .A3(new_n242_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1326gat));
  NAND3_X1  g442(.A1(new_n608_), .A2(new_n474_), .A3(new_n386_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n618_), .A2(new_n620_), .A3(new_n386_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(G22gat), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(G22gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT104), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n528_), .A2(new_n606_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n393_), .A2(new_n654_), .A3(new_n587_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n393_), .B2(new_n587_), .ZN(new_n657_));
  OAI211_X1 g456(.A(KEYINPUT44), .B(new_n653_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n652_), .B1(new_n659_), .B2(new_n655_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n661_));
  OAI211_X1 g460(.A(new_n658_), .B(new_n609_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G29gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n617_), .A2(new_n605_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n529_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n487_), .A3(new_n609_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT106), .ZN(G1328gat));
  NOR3_X1   g468(.A1(new_n665_), .A2(G36gat), .A3(new_n390_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G36gat), .B1(new_n673_), .B2(new_n390_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n672_), .A2(new_n674_), .A3(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  OAI21_X1  g478(.A(new_n493_), .B1(new_n665_), .B2(new_n638_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n242_), .A2(G43gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n673_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n666_), .B2(new_n386_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n673_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n385_), .A2(new_n491_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(G1331gat));
  NAND2_X1  g486(.A1(new_n607_), .A2(new_n472_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n689_), .A2(KEYINPUT108), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(KEYINPUT108), .ZN(new_n691_));
  AND4_X1   g490(.A1(new_n527_), .A2(new_n690_), .A3(new_n393_), .A4(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G57gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n609_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n618_), .A2(new_n605_), .A3(new_n527_), .A4(new_n472_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n380_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1332gat));
  INV_X1    g496(.A(G64gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(new_n698_), .A3(new_n631_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G64gat), .B1(new_n695_), .B2(new_n390_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT48), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n692_), .A2(new_n703_), .A3(new_n242_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G71gat), .B1(new_n695_), .B2(new_n638_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT49), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n692_), .A2(new_n708_), .A3(new_n386_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G78gat), .B1(new_n695_), .B2(new_n385_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1335gat));
  NAND4_X1  g512(.A1(new_n664_), .A2(new_n527_), .A3(new_n472_), .A4(new_n393_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT110), .ZN(new_n715_));
  AOI21_X1  g514(.A(G85gat), .B1(new_n715_), .B2(new_n609_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n472_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n527_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n717_), .A2(new_n605_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT111), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n609_), .A2(G85gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n716_), .B1(new_n721_), .B2(new_n722_), .ZN(G1336gat));
  AOI21_X1  g522(.A(G92gat), .B1(new_n715_), .B2(new_n631_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n631_), .A2(G92gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n721_), .B2(new_n725_), .ZN(G1337gat));
  NAND4_X1  g525(.A1(new_n715_), .A2(new_n400_), .A3(new_n402_), .A4(new_n242_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G99gat), .B1(new_n720_), .B2(new_n638_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT51), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1338gat));
  OAI211_X1 g532(.A(new_n386_), .B(new_n719_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT112), .B1(new_n734_), .B2(G106gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n738_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n385_), .A2(G106gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n715_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT53), .B1(new_n739_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n737_), .A2(new_n738_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n735_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n740_), .A4(new_n742_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(G1339gat));
  NAND2_X1  g548(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n602_), .A2(new_n604_), .A3(new_n527_), .A4(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n472_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n575_), .B(new_n752_), .C1(new_n586_), .C2(KEYINPUT37), .ZN(new_n753_));
  NOR2_X1   g552(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n562_), .A2(KEYINPUT76), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n579_), .A2(new_n576_), .A3(new_n546_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT77), .B1(new_n758_), .B2(new_n573_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n585_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n571_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n615_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n586_), .A2(KEYINPUT101), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n456_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT55), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n456_), .A2(new_n764_), .A3(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n442_), .A2(new_n455_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n766_), .B(new_n768_), .C1(new_n443_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(KEYINPUT56), .A4(new_n464_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n467_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n718_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n464_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n464_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(KEYINPUT115), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n774_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n523_), .B1(new_n506_), .B2(new_n518_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n517_), .B1(new_n516_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT116), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n525_), .A2(KEYINPUT117), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT117), .B1(new_n525_), .B2(new_n787_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n468_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n780_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n762_), .A2(new_n763_), .A3(KEYINPUT57), .A4(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n773_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n778_), .B2(new_n777_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n587_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n774_), .A2(new_n779_), .B1(new_n468_), .B2(new_n790_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n614_), .A2(new_n616_), .A3(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n793_), .B(new_n798_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n755_), .B1(new_n803_), .B2(new_n606_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n391_), .A2(new_n380_), .A3(new_n638_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n718_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n792_), .A2(KEYINPUT57), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n812_), .A2(new_n617_), .B1(new_n587_), .B2(new_n797_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n762_), .A2(new_n763_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n801_), .B1(new_n814_), .B2(new_n799_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n605_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT59), .B(new_n805_), .C1(new_n816_), .C2(new_n755_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n527_), .B1(new_n811_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n809_), .B1(new_n818_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n717_), .B2(KEYINPUT60), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n807_), .B(new_n821_), .C1(KEYINPUT60), .C2(new_n820_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n717_), .B1(new_n811_), .B2(new_n817_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n820_), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n807_), .A2(new_n825_), .A3(new_n605_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n606_), .B1(new_n811_), .B2(new_n817_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n825_), .ZN(G1342gat));
  INV_X1    g627(.A(G134gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n807_), .A2(new_n829_), .A3(new_n814_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n587_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n811_), .B2(new_n817_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(new_n829_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT120), .B(new_n830_), .C1(new_n832_), .C2(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1343gat));
  INV_X1    g636(.A(new_n804_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n385_), .A2(new_n242_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n390_), .A2(new_n839_), .A3(new_n609_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n718_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n472_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G148gat), .ZN(G1345gat));
  OAI211_X1 g644(.A(new_n605_), .B(new_n840_), .C1(new_n816_), .C2(new_n755_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  OR2_X1    g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n847_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1346gat));
  INV_X1    g652(.A(G162gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n841_), .A2(new_n854_), .A3(new_n814_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n841_), .A2(new_n587_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n854_), .ZN(G1347gat));
  NOR3_X1   g656(.A1(new_n390_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n838_), .A2(new_n718_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n859_), .A2(new_n860_), .A3(G169gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n838_), .A2(new_n858_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n718_), .A3(new_n300_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n859_), .B2(G169gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(G1348gat));
  AND3_X1   g665(.A1(new_n863_), .A2(G176gat), .A3(new_n472_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n472_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n215_), .B2(new_n868_), .ZN(G1349gat));
  NOR2_X1   g668(.A1(new_n862_), .A2(new_n606_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n870_), .B(new_n223_), .C1(new_n871_), .C2(G183gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT123), .A2(G183gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n870_), .B2(new_n873_), .ZN(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n862_), .B2(new_n831_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n814_), .A2(new_n224_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n862_), .B2(new_n876_), .ZN(G1351gat));
  NAND2_X1  g676(.A1(new_n839_), .A2(new_n380_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n631_), .B1(new_n878_), .B2(KEYINPUT124), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(KEYINPUT124), .B2(new_n878_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n838_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n883_));
  OR2_X1    g682(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n882_), .A2(new_n718_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n881_), .A2(new_n527_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n884_), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n472_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  AND2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n881_), .A2(new_n606_), .A3(new_n890_), .A4(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n882_), .A2(new_n605_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n890_), .ZN(G1354gat));
  NOR3_X1   g693(.A1(new_n881_), .A2(KEYINPUT126), .A3(new_n617_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(G218gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT126), .B1(new_n881_), .B2(new_n617_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n587_), .A2(G218gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT127), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n896_), .A2(new_n897_), .B1(new_n882_), .B2(new_n899_), .ZN(G1355gat));
endmodule


