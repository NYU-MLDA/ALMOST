//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  INV_X1    g002(.A(G71gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT77), .B(G43gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR3_X1   g007(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n209_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n218_), .A2(KEYINPUT75), .A3(KEYINPUT23), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT75), .B1(new_n218_), .B2(KEYINPUT23), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n218_), .B2(KEYINPUT23), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n218_), .A2(new_n229_), .A3(KEYINPUT23), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n221_), .A3(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n228_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT30), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G99gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT30), .B1(new_n225_), .B2(new_n236_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n208_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(new_n242_), .A3(new_n207_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n247_), .A3(KEYINPUT78), .ZN(new_n248_));
  INV_X1    g047(.A(G127gat), .ZN(new_n249_));
  INV_X1    g048(.A(G134gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G127gat), .A2(G134gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G113gat), .ZN(new_n254_));
  INV_X1    g053(.A(G113gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(G120gat), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(G120gat), .B1(new_n254_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT31), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(KEYINPUT31), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n248_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n245_), .A2(new_n247_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI211_X1 g067(.A(KEYINPUT78), .B(KEYINPUT79), .C1(new_n245_), .C2(new_n247_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n263_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n262_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  OR2_X1    g076(.A1(G211gat), .A2(G218gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G211gat), .A2(G218gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n276_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(KEYINPUT86), .A3(new_n279_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n277_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT87), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n277_), .A2(new_n284_), .A3(KEYINPUT87), .A4(new_n285_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n282_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(G141gat), .ZN(new_n292_));
  INV_X1    g091(.A(G148gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(G155gat), .A3(G162gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  INV_X1    g098(.A(G155gat), .ZN(new_n300_));
  INV_X1    g099(.A(G162gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT1), .B1(new_n300_), .B2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n291_), .B(new_n294_), .C1(new_n298_), .C2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n291_), .B1(new_n309_), .B2(KEYINPUT83), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT83), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n291_), .A2(KEYINPUT83), .A3(new_n309_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .A4(new_n316_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n302_), .A2(new_n303_), .B1(G155gat), .B2(G162gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n308_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n320_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(KEYINPUT2), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n313_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n314_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n308_), .B(new_n318_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n307_), .B1(new_n319_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n290_), .B1(new_n327_), .B2(KEYINPUT29), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(KEYINPUT88), .A2(G228gat), .A3(G233gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G78gat), .B(G106gat), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n332_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G22gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n319_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n325_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .A4(new_n307_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT28), .B1(new_n327_), .B2(KEYINPUT29), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n336_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n336_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(G50gat), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G50gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n343_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n346_), .A2(new_n349_), .A3(KEYINPUT85), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT85), .B1(new_n346_), .B2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n335_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n333_), .A2(KEYINPUT89), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n332_), .B(new_n353_), .Z(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n346_), .A3(new_n349_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G64gat), .ZN(new_n360_));
  INV_X1    g159(.A(G92gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n228_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n224_), .B2(new_n234_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT91), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT91), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n366_), .B(new_n363_), .C1(new_n224_), .C2(new_n234_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n231_), .A2(new_n221_), .A3(new_n232_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT90), .B1(new_n368_), .B2(new_n217_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n233_), .A2(new_n370_), .A3(new_n216_), .A4(new_n213_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n365_), .A2(new_n367_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n290_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n290_), .A2(new_n237_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n373_), .A2(KEYINPUT20), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n290_), .A2(new_n237_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT20), .B(new_n379_), .C1(new_n372_), .C2(new_n290_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n375_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n380_), .B2(new_n375_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n362_), .B(new_n378_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT100), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n233_), .A2(new_n216_), .A3(new_n213_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n290_), .A2(new_n386_), .A3(new_n364_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n237_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n375_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n375_), .B2(new_n380_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n362_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n384_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n380_), .A2(new_n375_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT92), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n380_), .A2(new_n381_), .A3(new_n375_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n397_), .A2(new_n385_), .A3(new_n362_), .A4(new_n378_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n357_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n391_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT27), .B1(new_n401_), .B2(new_n384_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n259_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n327_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n259_), .B(new_n307_), .C1(new_n319_), .C2(new_n326_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT94), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n405_), .A2(KEYINPUT4), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n405_), .A2(new_n412_), .A3(KEYINPUT4), .A4(new_n406_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n405_), .A2(new_n406_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n409_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT95), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT97), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT95), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n418_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n414_), .A2(new_n426_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n424_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n273_), .A2(new_n356_), .A3(new_n403_), .A4(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT101), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n429_), .A2(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT33), .B1(new_n436_), .B2(new_n425_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  NOR4_X1   g237(.A1(new_n429_), .A2(new_n430_), .A3(new_n438_), .A4(new_n424_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n408_), .A2(new_n409_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n415_), .A2(new_n410_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n424_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n362_), .B1(new_n397_), .B2(new_n378_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n384_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n401_), .A2(KEYINPUT93), .A3(new_n384_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n444_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n362_), .A2(KEYINPUT32), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT98), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n397_), .A3(new_n378_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n451_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n428_), .A2(new_n431_), .B1(new_n390_), .B2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n440_), .A2(new_n450_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n352_), .A2(new_n355_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT99), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n403_), .A2(new_n433_), .A3(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n390_), .A2(new_n454_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n432_), .A2(new_n453_), .A3(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n401_), .A2(KEYINPUT93), .A3(new_n384_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT93), .B1(new_n401_), .B2(new_n384_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n443_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n428_), .A2(new_n438_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n436_), .A2(KEYINPUT33), .A3(new_n425_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n461_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT99), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n356_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n458_), .A2(new_n459_), .A3(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n273_), .B(KEYINPUT80), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n435_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G127gat), .B(G155gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT16), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G183gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G211gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(G71gat), .B(G78gat), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(KEYINPUT11), .A3(new_n481_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G8gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n488_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT71), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n478_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT17), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n498_), .A2(new_n478_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT68), .B1(new_n511_), .B2(new_n506_), .ZN(new_n512_));
  INV_X1    g311(.A(G43gat), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n347_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n512_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G43gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n519_));
  AOI21_X1  g318(.A(G50gat), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n505_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n347_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(G50gat), .A3(new_n519_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT15), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n525_));
  INV_X1    g324(.A(G106gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n240_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT7), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT6), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n525_), .A2(new_n534_), .A3(new_n240_), .A4(new_n526_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n528_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G85gat), .B(G92gat), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n537_), .A2(KEYINPUT9), .B1(new_n530_), .B2(new_n532_), .ZN(new_n541_));
  INV_X1    g340(.A(G85gat), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n542_), .A2(new_n361_), .A3(KEYINPUT9), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT64), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT10), .B(G99gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(G106gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT10), .B(G99gat), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT64), .A3(new_n526_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n541_), .A2(new_n543_), .A3(new_n546_), .A4(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n536_), .A2(KEYINPUT8), .A3(new_n537_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n540_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n521_), .A2(new_n524_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n552_), .B(new_n554_), .C1(KEYINPUT35), .C2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n301_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT36), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n558_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n559_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n559_), .A2(new_n565_), .B1(new_n567_), .B2(new_n562_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT70), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT69), .B(new_n572_), .C1(new_n566_), .C2(new_n568_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(KEYINPUT37), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n573_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n474_), .A2(new_n504_), .A3(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n521_), .A2(new_n524_), .A3(new_n496_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT72), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT72), .B1(new_n522_), .B2(new_n523_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n495_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n521_), .A2(new_n586_), .A3(new_n524_), .A4(new_n496_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n580_), .A2(new_n581_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n581_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n584_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n496_), .B1(new_n590_), .B2(new_n582_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n583_), .A2(new_n584_), .A3(new_n495_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n227_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(G197gat), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n597_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(KEYINPUT74), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT74), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n594_), .A2(new_n602_), .A3(new_n597_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(G230gat), .ZN(new_n606_));
  INV_X1    g405(.A(G233gat), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n551_), .A2(new_n486_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n486_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n610_), .A2(new_n540_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(KEYINPUT12), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT12), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n551_), .A2(new_n613_), .A3(new_n486_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n608_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n608_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n618_), .B(new_n623_), .Z(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT67), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n578_), .A2(new_n605_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n490_), .A3(new_n432_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n474_), .A2(new_n604_), .A3(new_n627_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n569_), .B(KEYINPUT102), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n504_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n432_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G1gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n630_), .A2(new_n631_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n632_), .A2(KEYINPUT103), .A3(new_n639_), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1324gat));
  INV_X1    g444(.A(new_n403_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n629_), .A2(new_n491_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n637_), .A2(new_n646_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G8gat), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT39), .B(new_n491_), .C1(new_n637_), .C2(new_n646_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1325gat));
  NAND2_X1  g453(.A1(new_n637_), .A2(new_n472_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n655_), .B2(G15gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n629_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n473_), .A2(G15gat), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n656_), .A2(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(G1326gat));
  XNOR2_X1  g459(.A(new_n356_), .B(KEYINPUT104), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n629_), .A2(new_n336_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n637_), .A2(new_n661_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G22gat), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT42), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT42), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n503_), .A2(new_n569_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT106), .Z(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n633_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n432_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n448_), .A2(new_n449_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n465_), .A3(new_n466_), .A4(new_n443_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT99), .B(new_n457_), .C1(new_n675_), .C2(new_n461_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n469_), .B1(new_n468_), .B2(new_n356_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n472_), .B1(new_n678_), .B2(new_n459_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT43), .B(new_n577_), .C1(new_n679_), .C2(new_n435_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  INV_X1    g480(.A(new_n577_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n474_), .B2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n627_), .A2(new_n604_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n680_), .A2(new_n683_), .A3(new_n504_), .A4(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT105), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n685_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n433_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n673_), .B1(new_n690_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n689_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n646_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n403_), .B(KEYINPUT107), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n671_), .A2(new_n693_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n671_), .A2(KEYINPUT45), .A3(new_n693_), .A4(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n692_), .B1(new_n695_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n702_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n403_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n704_), .B(KEYINPUT46), .C1(new_n705_), .C2(new_n693_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1329gat));
  INV_X1    g506(.A(new_n689_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT44), .B1(new_n685_), .B2(KEYINPUT105), .ZN(new_n709_));
  OAI211_X1 g508(.A(G43gat), .B(new_n273_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n671_), .A2(new_n472_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT108), .B(G43gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n710_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  NAND3_X1  g517(.A1(new_n671_), .A2(new_n347_), .A3(new_n661_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n356_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n347_), .ZN(G1331gat));
  INV_X1    g520(.A(new_n627_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(new_n605_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n578_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n432_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n474_), .A2(new_n605_), .A3(new_n628_), .ZN(new_n726_));
  AND4_X1   g525(.A1(G57gat), .A2(new_n726_), .A3(new_n432_), .A4(new_n636_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1332gat));
  INV_X1    g527(.A(G64gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n729_), .A3(new_n697_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n726_), .A2(new_n636_), .A3(new_n697_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G64gat), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(KEYINPUT48), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(KEYINPUT48), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  NAND3_X1  g534(.A1(new_n724_), .A2(new_n204_), .A3(new_n472_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n726_), .A2(new_n636_), .A3(new_n472_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G71gat), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT49), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT49), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n724_), .A2(new_n742_), .A3(new_n661_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n636_), .A3(new_n661_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G78gat), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT50), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(KEYINPUT50), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n726_), .A2(new_n670_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n432_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n680_), .A2(new_n683_), .A3(new_n504_), .A4(new_n723_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n752_), .A2(new_n542_), .A3(new_n433_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1336gat));
  AOI21_X1  g553(.A(G92gat), .B1(new_n750_), .B2(new_n646_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n752_), .A2(new_n361_), .A3(new_n696_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1337gat));
  OAI21_X1  g556(.A(G99gat), .B1(new_n752_), .B2(new_n473_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(KEYINPUT109), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(G99gat), .C1(new_n752_), .C2(new_n473_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n273_), .A2(new_n547_), .ZN(new_n763_));
  OAI22_X1  g562(.A1(new_n759_), .A2(new_n762_), .B1(new_n749_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT51), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  OAI221_X1 g565(.A(new_n766_), .B1(new_n749_), .B2(new_n763_), .C1(new_n759_), .C2(new_n762_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1338gat));
  OAI21_X1  g567(.A(G106gat), .B1(new_n752_), .B2(new_n356_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT52), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(G106gat), .C1(new_n752_), .C2(new_n356_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n457_), .A2(new_n526_), .ZN(new_n774_));
  OAI22_X1  g573(.A1(new_n770_), .A2(new_n773_), .B1(new_n749_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  OAI221_X1 g576(.A(new_n777_), .B1(new_n749_), .B2(new_n774_), .C1(new_n770_), .C2(new_n773_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  NAND3_X1  g578(.A1(new_n612_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n615_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n615_), .A2(KEYINPUT111), .A3(KEYINPUT55), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT111), .B1(new_n615_), .B2(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n784_), .B(KEYINPUT112), .C1(new_n785_), .C2(new_n786_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n623_), .A3(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n618_), .A2(new_n623_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n601_), .A2(new_n603_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n789_), .A2(new_n623_), .A3(new_n790_), .A4(new_n792_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT114), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n580_), .A2(new_n589_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n581_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n597_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n600_), .A2(new_n803_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n624_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n794_), .A2(new_n797_), .A3(new_n806_), .A4(new_n798_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n569_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(KEYINPUT58), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n789_), .A2(new_n814_), .A3(new_n623_), .A4(new_n790_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n815_), .A2(new_n795_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n804_), .B1(new_n791_), .B2(KEYINPUT56), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n816_), .A2(new_n813_), .A3(new_n817_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n577_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n569_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n577_), .B(KEYINPUT116), .C1(new_n818_), .C2(new_n819_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n811_), .A2(new_n822_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n504_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n503_), .B(new_n604_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n827_), .B2(new_n627_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n576_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n504_), .B1(new_n829_), .B2(new_n574_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n604_), .A4(new_n722_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n834_), .ZN(new_n835_));
  AND4_X1   g634(.A1(new_n432_), .A2(new_n273_), .A3(new_n356_), .A4(new_n403_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n255_), .B1(new_n837_), .B2(new_n604_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT117), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n823_), .A2(new_n820_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n808_), .B2(new_n569_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n504_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT118), .B(new_n504_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n834_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n848_), .A2(new_n836_), .B1(KEYINPUT59), .B2(new_n837_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(G113gat), .A3(new_n605_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n839_), .A2(new_n850_), .ZN(G1340gat));
  INV_X1    g650(.A(new_n628_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n837_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n722_), .A2(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(KEYINPUT60), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(KEYINPUT60), .B2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n853_), .B2(new_n503_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n504_), .A2(new_n249_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n849_), .B2(new_n860_), .ZN(G1342gat));
  AOI21_X1  g660(.A(G134gat), .B1(new_n853_), .B2(new_n635_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n682_), .A2(new_n250_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n849_), .B2(new_n863_), .ZN(G1343gat));
  AOI21_X1  g663(.A(new_n833_), .B1(new_n825_), .B2(new_n504_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n472_), .A2(new_n356_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n697_), .A2(new_n433_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n865_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n605_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n852_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g673(.A1(new_n835_), .A2(new_n503_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT119), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n865_), .A2(new_n867_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n503_), .A4(new_n868_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n876_), .A2(new_n877_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n300_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n875_), .A2(KEYINPUT119), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n879_), .B1(new_n870_), .B2(new_n503_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT61), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n876_), .A2(new_n877_), .A3(new_n880_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G155gat), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n883_), .A2(new_n888_), .ZN(G1346gat));
  NAND3_X1  g688(.A1(new_n870_), .A2(G162gat), .A3(new_n577_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n870_), .A2(new_n635_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(G162gat), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1347gat));
  NAND3_X1  g693(.A1(new_n472_), .A2(new_n433_), .A3(new_n697_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n661_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n846_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT22), .B(G169gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n605_), .A2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT122), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT121), .B1(new_n897_), .B2(new_n604_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n846_), .A2(new_n904_), .A3(new_n605_), .A4(new_n896_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(G169gat), .A3(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n902_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n722_), .A2(G176gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n865_), .A2(new_n457_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n895_), .A2(new_n628_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n898_), .A2(new_n910_), .B1(new_n913_), .B2(G176gat), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT123), .Z(G1349gat));
  NOR3_X1   g714(.A1(new_n897_), .A2(new_n504_), .A3(new_n214_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n865_), .A2(new_n504_), .A3(new_n457_), .A4(new_n895_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT124), .ZN(new_n918_));
  INV_X1    g717(.A(G183gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n918_), .B2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n897_), .B2(new_n682_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n635_), .A2(new_n215_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n897_), .B2(new_n922_), .ZN(G1351gat));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n472_), .A2(new_n432_), .A3(new_n356_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n865_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n696_), .B1(new_n927_), .B2(KEYINPUT125), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n605_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n852_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g733(.A(KEYINPUT63), .B(G211gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n930_), .A2(new_n503_), .A3(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  OAI22_X1  g736(.A1(new_n929_), .A2(new_n504_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1354gat));
  OR3_X1    g740(.A1(new_n929_), .A2(KEYINPUT127), .A3(new_n634_), .ZN(new_n942_));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT127), .B1(new_n929_), .B2(new_n634_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n942_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n930_), .A2(G218gat), .A3(new_n577_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1355gat));
endmodule


