//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  XNOR2_X1  g000(.A(KEYINPUT79), .B(G15gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT78), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT23), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT75), .B(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n218_), .B2(G190gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n214_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(KEYINPUT25), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT25), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n207_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT24), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n216_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n227_), .A2(new_n231_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n220_), .A2(KEYINPUT30), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT30), .B1(new_n220_), .B2(new_n236_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n205_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n220_), .A2(new_n236_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT30), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n220_), .A2(new_n236_), .A3(KEYINPUT30), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n204_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  INV_X1    g044(.A(G43gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n239_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n203_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n244_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n239_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n202_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n255_), .A3(KEYINPUT81), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT31), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G113gat), .B(G120gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT80), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n250_), .A2(new_n255_), .A3(KEYINPUT81), .A4(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n257_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n257_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G22gat), .B(G50gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G228gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT85), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281_));
  INV_X1    g080(.A(G141gat), .ZN(new_n282_));
  INV_X1    g081(.A(G148gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n280_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n282_), .A2(new_n283_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(new_n285_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n279_), .B1(new_n277_), .B2(KEYINPUT1), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n300_));
  INV_X1    g099(.A(new_n279_), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n298_), .A2(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT82), .B(new_n279_), .C1(new_n277_), .C2(KEYINPUT1), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n297_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT29), .B1(new_n294_), .B2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT86), .B(G197gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(G204gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT21), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n313_));
  OR2_X1    g112(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n314_));
  INV_X1    g113(.A(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n310_), .B1(G197gat), .B2(G204gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n309_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n316_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(G204gat), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n306_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT21), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n312_), .B(new_n313_), .C1(new_n320_), .C2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n319_), .B(new_n309_), .C1(new_n308_), .C2(KEYINPUT21), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n313_), .B1(new_n328_), .B2(new_n312_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n276_), .B(new_n305_), .C1(new_n327_), .C2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n298_), .A2(new_n299_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n301_), .A2(new_n300_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n303_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n296_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n291_), .B(KEYINPUT83), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n279_), .B(new_n278_), .C1(new_n336_), .C2(new_n289_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n328_), .A2(new_n312_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n275_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n330_), .A2(G78gat), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(G78gat), .B1(new_n330_), .B2(new_n340_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n273_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n330_), .A2(new_n340_), .ZN(new_n344_));
  INV_X1    g143(.A(G78gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n330_), .A2(new_n340_), .A3(G78gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(G106gat), .A3(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n343_), .A2(new_n348_), .A3(KEYINPUT84), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT88), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n294_), .A2(new_n304_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n331_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT28), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n343_), .A2(new_n348_), .A3(KEYINPUT84), .A4(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n350_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n272_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n346_), .A2(new_n347_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n273_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n355_), .B1(new_n362_), .B2(new_n348_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n356_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n353_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n350_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n271_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n359_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT19), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n327_), .A2(new_n329_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n225_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT25), .B(G183gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n216_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n376_), .A2(new_n377_), .B1(new_n212_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n328_), .A2(new_n312_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n240_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n371_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n379_), .A2(new_n339_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n339_), .A2(new_n236_), .A3(new_n220_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n385_), .A2(KEYINPUT20), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n387_), .B2(new_n371_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n385_), .A2(KEYINPUT20), .A3(new_n370_), .A4(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n379_), .A2(new_n339_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n370_), .B1(new_n383_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT93), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n388_), .B(new_n394_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n393_), .B1(new_n399_), .B2(KEYINPUT93), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n264_), .A2(new_n351_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n351_), .A2(new_n260_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n264_), .A2(new_n351_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(KEYINPUT4), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  AOI21_X1  g213(.A(new_n408_), .B1(new_n351_), .B2(new_n260_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n407_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n410_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n414_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n401_), .A2(new_n402_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n392_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n383_), .A2(new_n397_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n371_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n392_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n395_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT90), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT33), .B(new_n414_), .C1(new_n410_), .C2(new_n417_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n407_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n427_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT91), .B(KEYINPUT33), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n419_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT92), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT92), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n419_), .A2(new_n440_), .A3(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n420_), .B1(new_n435_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n270_), .B1(new_n368_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n424_), .B1(new_n423_), .B2(new_n395_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n388_), .A2(new_n392_), .B1(new_n445_), .B2(KEYINPUT94), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n445_), .A2(KEYINPUT94), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT27), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n426_), .A2(KEYINPUT27), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n418_), .A2(new_n419_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n359_), .A2(new_n453_), .A3(new_n367_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n450_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n359_), .B2(new_n367_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n268_), .A2(new_n269_), .A3(new_n451_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n444_), .A2(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  INV_X1    g258(.A(G1gat), .ZN(new_n460_));
  INV_X1    g259(.A(G8gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G8gat), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n464_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n470_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(KEYINPUT15), .A3(new_n470_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n467_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT73), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n485_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT74), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n458_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n494_));
  INV_X1    g293(.A(G85gat), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n493_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT9), .A3(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n273_), .A3(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n498_), .A2(new_n503_), .A3(new_n506_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n505_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n515_), .B2(new_n503_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n510_), .B1(new_n516_), .B2(KEYINPUT8), .ZN(new_n517_));
  INV_X1    g316(.A(new_n511_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT8), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520_));
  INV_X1    g319(.A(G99gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n273_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n512_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n523_), .A2(KEYINPUT65), .B1(new_n500_), .B2(new_n502_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(new_n525_), .A3(new_n512_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n492_), .B1(new_n517_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(KEYINPUT65), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n526_), .A3(new_n503_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n519_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n503_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n518_), .B1(new_n533_), .B2(new_n523_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n532_), .A2(new_n536_), .A3(KEYINPUT67), .A4(new_n510_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n528_), .A2(new_n537_), .A3(new_n481_), .A4(new_n480_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT70), .B1(new_n540_), .B2(KEYINPUT35), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n517_), .A2(new_n527_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n473_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(KEYINPUT35), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n538_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  OR4_X1    g348(.A1(KEYINPUT36), .A2(new_n545_), .A3(new_n546_), .A4(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(KEYINPUT36), .Z(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n553_), .A2(KEYINPUT37), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(KEYINPUT37), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n467_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(G64gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(G57gat), .ZN(new_n565_));
  INV_X1    g364(.A(G57gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(G64gat), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n565_), .A2(new_n567_), .A3(KEYINPUT66), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT66), .B1(new_n565_), .B2(new_n567_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT11), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT66), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT11), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n567_), .A3(KEYINPUT66), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G71gat), .B(G78gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT11), .B(new_n577_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n563_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n561_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n561_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT17), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n557_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n542_), .A2(new_n581_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n542_), .A2(new_n581_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n579_), .A2(KEYINPUT12), .A3(new_n580_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n528_), .A3(new_n537_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n542_), .B2(new_n581_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n593_), .B1(new_n542_), .B2(new_n581_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G120gat), .B(G148gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT5), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT68), .B1(new_n603_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n596_), .A2(new_n602_), .A3(new_n610_), .A4(new_n607_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n609_), .A2(new_n611_), .B1(new_n603_), .B2(new_n608_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT69), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT13), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT13), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n592_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n491_), .A2(KEYINPUT95), .A3(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n357_), .A2(new_n358_), .A3(new_n272_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n271_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n443_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n270_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n454_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n456_), .A2(new_n457_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n490_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n619_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n620_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n460_), .A3(new_n451_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n627_), .A2(new_n553_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(KEYINPUT96), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(KEYINPUT96), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n489_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n618_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n591_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n460_), .B1(new_n643_), .B2(new_n451_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n635_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  NOR2_X1   g445(.A1(new_n450_), .A2(G8gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n620_), .A2(new_n631_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n642_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n455_), .B(new_n651_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n461_), .B1(new_n653_), .B2(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(KEYINPUT39), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n652_), .B(new_n654_), .C1(new_n653_), .C2(KEYINPUT39), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n650_), .A2(new_n657_), .A3(new_n658_), .A4(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OAI211_X1 g463(.A(new_n270_), .B(new_n651_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G15gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT41), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n668_), .A3(G15gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n667_), .A2(KEYINPUT100), .A3(new_n669_), .ZN(new_n673_));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n632_), .A2(new_n674_), .A3(new_n270_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT101), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n673_), .A3(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n368_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n632_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n643_), .A2(new_n679_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G22gat), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT42), .B(new_n678_), .C1(new_n643_), .C2(new_n679_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1327gat));
  INV_X1    g484(.A(new_n591_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n553_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n618_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n491_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n451_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n458_), .B2(new_n557_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n627_), .A2(KEYINPUT43), .A3(new_n556_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(new_n686_), .A3(new_n641_), .A4(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n627_), .A2(new_n556_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n591_), .B1(new_n699_), .B2(new_n693_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n641_), .A4(new_n695_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n451_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n692_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  XOR2_X1   g503(.A(new_n450_), .B(KEYINPUT102), .Z(new_n705_));
  NOR3_X1   g504(.A1(new_n690_), .A2(G36gat), .A3(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n698_), .A2(new_n701_), .A3(new_n455_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(KEYINPUT46), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1329gat));
  XNOR2_X1  g514(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n624_), .A2(new_n246_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n698_), .A2(new_n701_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n246_), .B1(new_n690_), .B2(new_n624_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n716_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1330gat));
  AOI21_X1  g528(.A(G50gat), .B1(new_n691_), .B2(new_n679_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n679_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n702_), .B2(new_n731_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n592_), .A2(new_n617_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT106), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(new_n458_), .A3(new_n489_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n451_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT107), .Z(new_n737_));
  NOR4_X1   g536(.A1(new_n639_), .A2(new_n628_), .A3(new_n617_), .A4(new_n686_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n452_), .A2(new_n566_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(G1332gat));
  INV_X1    g539(.A(new_n705_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n564_), .A3(new_n741_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n686_), .A2(new_n628_), .A3(new_n617_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n741_), .B(new_n743_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G64gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT109), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n747_), .A3(G64gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n746_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n742_), .B1(new_n750_), .B2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n735_), .A2(new_n753_), .A3(new_n270_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n270_), .B(new_n743_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G71gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT111), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n758_), .A3(G71gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n760_));
  AND3_X1   g559(.A1(new_n757_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n754_), .B1(new_n761_), .B2(new_n762_), .ZN(G1334gat));
  NAND3_X1  g562(.A1(new_n735_), .A2(new_n345_), .A3(new_n679_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n679_), .B(new_n743_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G78gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G78gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT112), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n764_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1335gat));
  NOR4_X1   g572(.A1(new_n458_), .A2(new_n489_), .A3(new_n617_), .A4(new_n688_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n451_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT113), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n617_), .A2(new_n489_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n700_), .A2(new_n695_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n451_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n776_), .A2(new_n780_), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n778_), .B2(new_n705_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n774_), .A2(new_n493_), .A3(new_n455_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n778_), .B2(new_n624_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n270_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n774_), .A2(new_n786_), .B1(KEYINPUT114), .B2(KEYINPUT51), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n788_), .B(new_n789_), .Z(G1338gat));
  NAND3_X1  g589(.A1(new_n774_), .A2(new_n273_), .A3(new_n679_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n700_), .A2(new_n679_), .A3(new_n695_), .A4(new_n777_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n792_), .B2(G106gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n791_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n557_), .A2(new_n490_), .A3(new_n591_), .A4(new_n617_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n609_), .A2(new_n611_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(new_n489_), .A3(KEYINPUT115), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT115), .B1(new_n806_), .B2(new_n489_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n602_), .A2(KEYINPUT55), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n598_), .A2(new_n600_), .A3(new_n601_), .A4(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n542_), .A2(new_n581_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n598_), .A2(new_n600_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n593_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(KEYINPUT116), .A3(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n608_), .ZN(new_n822_));
  AOI221_X4 g621(.A(new_n818_), .B1(new_n815_), .B2(new_n593_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n813_), .B2(new_n816_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT56), .B(new_n608_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n809_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n484_), .A2(new_n488_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n475_), .A2(new_n476_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n482_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n488_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n612_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n687_), .B1(new_n827_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n608_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n825_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n832_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n841_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n839_), .B2(new_n825_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT58), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n556_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n833_), .B1(new_n840_), .B2(new_n809_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n687_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n836_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n805_), .B1(new_n686_), .B2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n624_), .A2(new_n452_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n456_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n802_), .B1(new_n857_), .B2(new_n640_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(KEYINPUT117), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n556_), .B1(new_n846_), .B2(KEYINPUT58), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n843_), .B(new_n845_), .C1(new_n839_), .C2(new_n825_), .ZN(new_n861_));
  OAI22_X1  g660(.A1(new_n835_), .A2(KEYINPUT57), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n848_), .A2(new_n864_), .A3(new_n851_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n836_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n805_), .B1(new_n866_), .B2(new_n686_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n854_), .A2(new_n456_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n857_), .B2(KEYINPUT59), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT120), .B(G113gat), .Z(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n628_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n858_), .A2(KEYINPUT117), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n859_), .A2(new_n873_), .A3(new_n874_), .ZN(G1340gat));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n617_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n856_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n871_), .A2(new_n618_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n876_), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n871_), .A2(G127gat), .A3(new_n591_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G127gat), .B1(new_n856_), .B2(new_n591_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n884_), .A3(new_n885_), .ZN(G1342gat));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n853_), .B2(new_n855_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n887_), .B(new_n556_), .C1(new_n867_), .C2(new_n869_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G134gat), .ZN(new_n889_));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n856_), .A2(new_n890_), .A3(new_n687_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n889_), .A2(KEYINPUT122), .A3(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1343gat));
  NOR2_X1   g695(.A1(new_n853_), .A2(new_n368_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n897_), .A2(new_n451_), .A3(new_n624_), .A4(new_n705_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n640_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n282_), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n617_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n283_), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n898_), .A2(new_n686_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n898_), .B2(new_n557_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n553_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n898_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  INV_X1    g708(.A(new_n457_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n705_), .A2(new_n910_), .A3(new_n679_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n867_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n489_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n909_), .B1(new_n914_), .B2(G169gat), .ZN(new_n915_));
  AOI211_X1 g714(.A(KEYINPUT62), .B(new_n228_), .C1(new_n913_), .C2(new_n489_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n867_), .B2(new_n912_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n862_), .A2(KEYINPUT119), .B1(KEYINPUT57), .B2(new_n835_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n591_), .B1(new_n919_), .B2(new_n865_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n911_), .B(KEYINPUT123), .C1(new_n920_), .C2(new_n805_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n489_), .A2(new_n206_), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT124), .Z(new_n925_));
  OAI22_X1  g724(.A1(new_n915_), .A2(new_n916_), .B1(new_n923_), .B2(new_n925_), .ZN(G1348gat));
  NOR2_X1   g725(.A1(new_n853_), .A2(new_n912_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(G176gat), .A3(new_n618_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n617_), .B1(new_n918_), .B2(new_n921_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(G176gat), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(KEYINPUT125), .B(new_n928_), .C1(new_n929_), .C2(G176gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1349gat));
  AOI21_X1  g733(.A(new_n218_), .B1(new_n927_), .B2(new_n591_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n686_), .A2(new_n375_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n922_), .B2(new_n936_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n923_), .B2(new_n557_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n922_), .A2(new_n374_), .A3(new_n687_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1351gat));
  NAND4_X1  g739(.A1(new_n897_), .A2(new_n452_), .A3(new_n624_), .A4(new_n741_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n640_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT126), .B(G197gat), .Z(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1352gat));
  NOR2_X1   g743(.A1(new_n941_), .A2(new_n617_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n945_), .B1(KEYINPUT127), .B2(new_n315_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT127), .B(G204gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n945_), .B2(new_n947_), .ZN(G1353gat));
  NOR2_X1   g747(.A1(new_n941_), .A2(new_n686_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  AND2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n949_), .B2(new_n950_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n941_), .B2(new_n557_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n553_), .A2(G218gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n941_), .B2(new_n955_), .ZN(G1355gat));
endmodule


