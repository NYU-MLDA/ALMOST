//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n594_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT71), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT70), .B(G15gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(G22gat), .ZN(new_n212_));
  INV_X1    g011(.A(G1gat), .ZN(new_n213_));
  INV_X1    g012(.A(G8gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G1gat), .B(G8gat), .Z(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n217_), .A3(new_n215_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n210_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n220_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT72), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n221_), .B(new_n222_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n208_), .B(KEYINPUT71), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n222_), .B1(new_n230_), .B2(new_n221_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G169gat), .B(G197gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(KEYINPUT73), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n233_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  INV_X1    g039(.A(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(G15gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n242_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G169gat), .ZN(new_n246_));
  INV_X1    g045(.A(G176gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT24), .ZN(new_n258_));
  INV_X1    g057(.A(G169gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n247_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n254_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n251_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n262_), .B(new_n265_), .C1(new_n258_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT76), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT76), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n245_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n245_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G113gat), .B(G120gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT77), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n279_), .B(KEYINPUT31), .Z(new_n280_));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n280_), .A2(new_n281_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n273_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT3), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(KEYINPUT3), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n294_), .A2(new_n297_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n290_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n289_), .B(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n293_), .B(new_n295_), .C1(new_n303_), .C2(new_n288_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n279_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n304_), .A3(new_n277_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(KEYINPUT4), .A3(new_n307_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n309_), .B(KEYINPUT92), .Z(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n313_));
  NAND3_X1  g112(.A1(new_n279_), .A2(new_n305_), .A3(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G29gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G85gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT0), .B(G57gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n310_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n284_), .B1(new_n273_), .B2(new_n283_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n285_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT86), .ZN(new_n334_));
  XOR2_X1   g133(.A(G211gat), .B(G218gat), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(KEYINPUT86), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(KEYINPUT21), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G204gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT83), .A3(G197gat), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT21), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n337_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n346_), .A3(new_n339_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(KEYINPUT87), .A3(new_n337_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n268_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n254_), .B1(new_n261_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n357_), .B(new_n265_), .C1(new_n266_), .C2(new_n356_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n248_), .A2(new_n251_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n256_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n349_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT20), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n332_), .B1(new_n355_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT91), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NOR2_X1   g168(.A1(new_n361_), .A2(new_n349_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n351_), .A2(new_n268_), .A3(new_n354_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n331_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n375_), .B(new_n332_), .C1(new_n355_), .C2(new_n363_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n365_), .A2(new_n369_), .A3(new_n374_), .A4(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n377_), .A2(KEYINPUT27), .ZN(new_n378_));
  INV_X1    g177(.A(new_n369_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n331_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT95), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n257_), .A2(new_n267_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n349_), .A2(new_n350_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT87), .B1(new_n353_), .B2(new_n337_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n371_), .B1(new_n361_), .B2(new_n349_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n380_), .A2(new_n381_), .B1(new_n387_), .B2(new_n332_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n380_), .A2(new_n381_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n379_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n376_), .A2(new_n374_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n375_), .B1(new_n387_), .B2(new_n332_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n379_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n377_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n378_), .A2(new_n390_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT80), .B(KEYINPUT28), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G22gat), .B(G50gat), .Z(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  AND2_X1   g200(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(G228gat), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT82), .Z(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n305_), .B2(KEYINPUT29), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT88), .ZN(new_n408_));
  XOR2_X1   g207(.A(G78gat), .B(G106gat), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n404_), .B1(new_n411_), .B2(new_n349_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n407_), .B2(KEYINPUT88), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n401_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n399_), .B(new_n400_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n414_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT96), .B1(new_n396_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n394_), .A2(new_n395_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n390_), .A2(KEYINPUT27), .A3(new_n377_), .ZN(new_n424_));
  AND4_X1   g223(.A1(KEYINPUT96), .A2(new_n423_), .A3(new_n424_), .A4(new_n421_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n328_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n285_), .A2(new_n326_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n417_), .A2(new_n420_), .ZN(new_n428_));
  AND4_X1   g227(.A1(new_n428_), .A2(new_n325_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n365_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n431_), .B(new_n324_), .C1(new_n430_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(KEYINPUT33), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n310_), .A2(new_n315_), .A3(new_n320_), .A4(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n308_), .A2(new_n312_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n311_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n321_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n323_), .A2(new_n435_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n393_), .A3(new_n377_), .A4(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n428_), .B1(new_n433_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n427_), .B1(new_n429_), .B2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n239_), .B1(new_n426_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G232gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT34), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT35), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT68), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT69), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT10), .B(G99gat), .Z(new_n453_));
  AND2_X1   g252(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT6), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n459_), .A2(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n466_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n459_), .A2(new_n461_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473_));
  INV_X1    g272(.A(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT7), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n469_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n468_), .B1(new_n478_), .B2(KEYINPUT8), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n459_), .A2(new_n461_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n473_), .A2(new_n471_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n466_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT8), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n452_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n453_), .A2(new_n456_), .B1(new_n466_), .B2(KEYINPUT9), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n483_), .A2(new_n484_), .B1(new_n464_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n478_), .A2(KEYINPUT8), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT66), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n208_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n448_), .A2(KEYINPUT35), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n489_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n225_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n451_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n450_), .A2(KEYINPUT69), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n491_), .A2(new_n494_), .A3(KEYINPUT69), .A4(new_n450_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G190gat), .B(G218gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(KEYINPUT36), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n503_), .B(KEYINPUT36), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n498_), .A2(new_n499_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT37), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n479_), .A2(new_n485_), .A3(new_n452_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT66), .B1(new_n488_), .B2(new_n489_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n522_));
  INV_X1    g321(.A(new_n518_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n486_), .A2(new_n523_), .A3(new_n490_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n486_), .A2(new_n490_), .A3(KEYINPUT67), .A4(new_n523_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n493_), .A2(KEYINPUT12), .A3(new_n518_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n521_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n533_), .A3(new_n526_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT5), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n529_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n511_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n529_), .A2(new_n534_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n538_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n529_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT13), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n223_), .A2(new_n518_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n523_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT16), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n552_), .A2(KEYINPUT17), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n556_), .B(KEYINPUT17), .ZN(new_n560_));
  INV_X1    g359(.A(new_n558_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n560_), .B1(new_n561_), .B2(new_n551_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n510_), .A2(new_n547_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n446_), .A2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n565_), .A2(G1gat), .A3(new_n325_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT97), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT38), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT38), .ZN(new_n569_));
  INV_X1    g368(.A(new_n508_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n426_), .B2(new_n445_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n547_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n238_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n563_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G1gat), .B1(new_n575_), .B2(new_n325_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n569_), .A3(new_n576_), .ZN(G1324gat));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n396_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n214_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n446_), .A2(new_n214_), .A3(new_n579_), .A4(new_n564_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(G1325gat));
  OAI21_X1  g385(.A(G15gat), .B1(new_n575_), .B2(new_n427_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT41), .Z(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT100), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT100), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n565_), .A2(G15gat), .A3(new_n427_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT101), .Z(new_n592_));
  NAND3_X1  g391(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(G1326gat));
  OAI21_X1  g392(.A(G22gat), .B1(new_n575_), .B2(new_n421_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT42), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n421_), .A2(G22gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n565_), .B2(new_n596_), .ZN(G1327gat));
  NAND2_X1  g396(.A1(new_n570_), .A2(new_n563_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n547_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n446_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G29gat), .B1(new_n601_), .B2(new_n324_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n396_), .A2(KEYINPUT96), .A3(new_n421_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n423_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n327_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n427_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n433_), .A2(new_n443_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n421_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n428_), .A2(new_n325_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n510_), .B(new_n603_), .C1(new_n608_), .C2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n509_), .B1(new_n426_), .B2(new_n445_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n563_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n573_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT102), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT104), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n623_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n625_), .A3(new_n620_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n324_), .A2(G29gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n602_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  INV_X1    g428(.A(KEYINPUT106), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT46), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(KEYINPUT46), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n396_), .A2(G36gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n600_), .A2(KEYINPUT45), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT45), .B1(new_n600_), .B2(new_n634_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n617_), .A2(new_n625_), .A3(new_n620_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n625_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT105), .B(new_n579_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G36gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT105), .B1(new_n627_), .B2(new_n579_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n631_), .B(new_n637_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n579_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(G36gat), .A3(new_n640_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n631_), .B1(new_n648_), .B2(new_n637_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n644_), .A2(new_n649_), .ZN(G1329gat));
  XOR2_X1   g449(.A(KEYINPUT107), .B(G43gat), .Z(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n601_), .B2(new_n609_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n427_), .A2(new_n241_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n627_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g454(.A1(new_n421_), .A2(G50gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT108), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n601_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n421_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n659_));
  INV_X1    g458(.A(G50gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT109), .ZN(G1331gat));
  NOR2_X1   g461(.A1(new_n233_), .A2(new_n237_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n237_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n663_), .A2(new_n563_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n571_), .A2(new_n547_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G57gat), .B1(new_n667_), .B2(new_n325_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n238_), .B1(new_n426_), .B2(new_n445_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n669_), .A2(new_n547_), .A3(new_n618_), .A4(new_n509_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n325_), .A2(G57gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1332gat));
  OAI21_X1  g471(.A(G64gat), .B1(new_n667_), .B2(new_n396_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT48), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n396_), .A2(G64gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n670_), .B2(new_n675_), .ZN(G1333gat));
  OAI21_X1  g475(.A(G71gat), .B1(new_n667_), .B2(new_n427_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT49), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n427_), .A2(G71gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n670_), .B2(new_n679_), .ZN(G1334gat));
  OAI21_X1  g479(.A(G78gat), .B1(new_n667_), .B2(new_n421_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT50), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n421_), .A2(G78gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n670_), .B2(new_n683_), .ZN(G1335gat));
  NOR3_X1   g483(.A1(new_n572_), .A2(new_n238_), .A3(new_n618_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n617_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n510_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n616_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT110), .A3(new_n614_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n686_), .B1(new_n688_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G85gat), .B1(new_n694_), .B2(new_n325_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n572_), .A2(new_n598_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n669_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G85gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n324_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n697_), .B2(new_n699_), .ZN(G1336gat));
  OAI21_X1  g499(.A(G92gat), .B1(new_n694_), .B2(new_n396_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n697_), .A2(G92gat), .A3(new_n396_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1337gat));
  NAND2_X1  g505(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n609_), .A2(new_n453_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n697_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n693_), .A2(new_n609_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G99gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(G1338gat));
  NAND4_X1  g512(.A1(new_n669_), .A2(new_n428_), .A3(new_n456_), .A4(new_n696_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n685_), .A2(new_n428_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n691_), .B2(new_n614_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(G106gat), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT113), .B1(new_n716_), .B2(new_n475_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n714_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT53), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n714_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1339gat));
  AOI211_X1 g527(.A(new_n325_), .B(new_n427_), .C1(new_n604_), .C2(new_n607_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n236_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n222_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n221_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n223_), .A2(new_n225_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT72), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n733_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n732_), .B1(new_n230_), .B2(new_n221_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n731_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n222_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n236_), .B1(new_n741_), .B2(new_n231_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n739_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n545_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n523_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n530_), .B(new_n524_), .C1(new_n748_), .C2(KEYINPUT12), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(new_n527_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n527_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n531_), .A2(new_n533_), .A3(KEYINPUT55), .A4(new_n526_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n538_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n526_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n534_), .B1(new_n758_), .B2(new_n747_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n753_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n538_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n746_), .B1(new_n757_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT58), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n745_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n739_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n540_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n538_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n756_), .B(new_n539_), .C1(new_n759_), .C2(new_n753_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(KEYINPUT117), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n510_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n238_), .A2(new_n545_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n765_), .A2(new_n766_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n508_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n774_), .B1(new_n757_), .B2(new_n761_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n508_), .B1(new_n783_), .B2(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n780_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n773_), .A2(new_n782_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n563_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n542_), .A2(new_n546_), .A3(new_n666_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n542_), .A2(new_n546_), .A3(new_n666_), .A4(KEYINPUT114), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n509_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT54), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n790_), .A2(new_n794_), .A3(new_n509_), .A4(new_n791_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n730_), .B1(new_n787_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(G113gat), .B1(new_n798_), .B2(new_n238_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT59), .B1(new_n798_), .B2(KEYINPUT118), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n796_), .B1(new_n786_), .B2(new_n563_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .A4(new_n730_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT119), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n781_), .B1(new_n779_), .B2(new_n508_), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n570_), .B(new_n780_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n618_), .B1(new_n808_), .B2(new_n773_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT118), .B(new_n729_), .C1(new_n809_), .C2(new_n796_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n803_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n798_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n805_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n238_), .A2(G113gat), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT120), .Z(new_n817_));
  AOI21_X1  g616(.A(new_n799_), .B1(new_n815_), .B2(new_n817_), .ZN(G1340gat));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n572_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n798_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT121), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n572_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n819_), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n563_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n805_), .A2(new_n814_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n798_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n828_), .B2(new_n563_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(KEYINPUT122), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1342gat));
  NAND3_X1  g633(.A1(new_n805_), .A2(new_n814_), .A3(new_n510_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G134gat), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n508_), .A2(G134gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n828_), .B2(new_n837_), .ZN(G1343gat));
  NOR3_X1   g637(.A1(new_n801_), .A2(new_n421_), .A3(new_n609_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n579_), .A2(new_n325_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n239_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT123), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n572_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n292_), .ZN(G1345gat));
  AND2_X1   g645(.A1(new_n839_), .A2(new_n840_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n618_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT124), .B1(new_n841_), .B2(new_n563_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n851_), .B(new_n853_), .ZN(G1346gat));
  OR3_X1    g653(.A1(new_n841_), .A2(G162gat), .A3(new_n508_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G162gat), .B1(new_n841_), .B2(new_n509_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n787_), .A2(new_n797_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n327_), .A2(new_n396_), .A3(new_n428_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n238_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT125), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n259_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n858_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n858_), .A3(new_n865_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(KEYINPUT62), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n866_), .A2(new_n870_), .B1(new_n246_), .B2(new_n862_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1348gat));
  NAND2_X1  g671(.A1(new_n859_), .A2(new_n860_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n572_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n247_), .ZN(G1349gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n563_), .ZN(new_n876_));
  MUX2_X1   g675(.A(G183gat), .B(new_n263_), .S(new_n876_), .Z(G1350gat));
  OAI21_X1  g676(.A(G190gat), .B1(new_n873_), .B2(new_n509_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n570_), .A2(new_n264_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n873_), .B2(new_n879_), .ZN(G1351gat));
  NOR2_X1   g679(.A1(new_n396_), .A2(new_n324_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n839_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n238_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n572_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n342_), .ZN(G1353gat));
  NOR2_X1   g686(.A1(new_n882_), .A2(new_n563_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  AND2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n888_), .B2(new_n889_), .ZN(G1354gat));
  AOI21_X1  g691(.A(G218gat), .B1(new_n883_), .B2(new_n570_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n510_), .A2(G218gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT127), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n883_), .B2(new_n895_), .ZN(G1355gat));
endmodule


