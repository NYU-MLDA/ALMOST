//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n203_), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n208_), .B(new_n209_), .C1(new_n210_), .C2(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n212_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n203_), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT66), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n207_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT8), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n211_), .A2(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n219_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT64), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(KEYINPUT64), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT10), .B(G99gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n209_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n215_), .A2(new_n216_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n225_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(new_n224_), .A3(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G57gat), .B(G64gat), .Z(new_n235_));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n239_));
  XOR2_X1   g038(.A(G71gat), .B(G78gat), .Z(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n239_), .A2(new_n240_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n234_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n243_), .A2(new_n220_), .A3(new_n224_), .A4(new_n233_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n234_), .A2(new_n248_), .A3(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n246_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT67), .B(G204gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G120gat), .B(G148gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT5), .B(G176gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n252_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT13), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT13), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G8gat), .B(G36gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT87), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT19), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT85), .B(G197gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT21), .B(new_n281_), .C1(new_n282_), .C2(G204gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G197gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n283_), .B(new_n285_), .C1(new_n288_), .C2(KEYINPUT21), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n284_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT80), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(G183gat), .A3(G190gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n293_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n294_), .A2(new_n296_), .A3(KEYINPUT81), .A4(new_n297_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT24), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  MUX2_X1   g106(.A(new_n306_), .B(KEYINPUT24), .S(new_n307_), .Z(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT26), .B(G190gat), .Z(new_n309_));
  OR2_X1    g108(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n304_), .B(new_n308_), .C1(new_n309_), .C2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n301_), .A2(new_n293_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n297_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G183gat), .ZN(new_n317_));
  INV_X1    g116(.A(G190gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n305_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n292_), .B1(new_n313_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n308_), .B1(new_n315_), .B2(new_n314_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n310_), .A2(KEYINPUT89), .A3(new_n311_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT89), .B1(new_n310_), .B2(new_n311_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n309_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n324_), .B1(new_n304_), .B2(new_n319_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n334_), .A2(new_n291_), .A3(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n327_), .B1(new_n339_), .B2(KEYINPUT98), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n280_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n292_), .A2(new_n326_), .A3(new_n313_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT90), .B1(new_n328_), .B2(new_n333_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n346_));
  INV_X1    g145(.A(new_n309_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n316_), .A2(new_n346_), .A3(new_n308_), .A4(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n335_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT20), .B(new_n344_), .C1(new_n350_), .C2(new_n292_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n279_), .B(KEYINPUT88), .Z(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n276_), .B1(new_n343_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT84), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT2), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G141gat), .A2(G148gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(KEYINPUT84), .A3(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n361_), .A2(new_n364_), .A3(new_n365_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT1), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n358_), .A2(new_n369_), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n362_), .B1(new_n356_), .B2(KEYINPUT1), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n358_), .A2(new_n368_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G113gat), .ZN(new_n375_));
  INV_X1    g174(.A(G134gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G113gat), .A2(G134gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G120gat), .ZN(new_n380_));
  INV_X1    g179(.A(G120gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n380_), .A2(G127gat), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(G127gat), .B1(new_n380_), .B2(new_n382_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(new_n384_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n373_), .A3(new_n372_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n388_), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n387_), .A2(new_n372_), .A3(KEYINPUT4), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n355_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G85gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(G1gat), .B(G29gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n355_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n397_));
  OR3_X1    g196(.A1(new_n391_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n391_), .B2(new_n397_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT99), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT99), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(new_n395_), .C1(new_n391_), .C2(new_n397_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n351_), .A2(new_n352_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n345_), .A2(new_n349_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n335_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n292_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n327_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n350_), .A2(KEYINPUT91), .A3(new_n292_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n408_), .A2(KEYINPUT20), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n275_), .B(new_n403_), .C1(new_n411_), .C2(new_n279_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n354_), .A2(new_n400_), .A3(new_n402_), .A4(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n403_), .B1(new_n411_), .B2(new_n279_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n274_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n274_), .B(new_n403_), .C1(new_n411_), .C2(new_n279_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n389_), .A2(new_n390_), .A3(new_n355_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n395_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n386_), .A2(new_n388_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT95), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n386_), .A2(KEYINPUT95), .A3(new_n388_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n396_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT96), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n420_), .A2(new_n428_), .A3(new_n425_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n416_), .A2(new_n417_), .A3(new_n427_), .A4(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n399_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n413_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n372_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n291_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n438_), .A2(G228gat), .A3(G233gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(G228gat), .B2(G233gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n372_), .A2(new_n436_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G22gat), .B(G50gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT28), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n444_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G78gat), .B(G106gat), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n445_), .B(new_n446_), .C1(KEYINPUT86), .C2(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n441_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n451_), .B(new_n450_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT30), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT31), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n458_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n387_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n458_), .B(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n385_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G99gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n326_), .A2(new_n469_), .A3(new_n313_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n326_), .B2(new_n313_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n326_), .A2(new_n313_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT82), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(KEYINPUT83), .A3(new_n470_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n467_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(new_n476_), .A3(new_n467_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n465_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n473_), .A2(new_n476_), .A3(new_n467_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n462_), .A2(new_n464_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n435_), .A2(new_n455_), .A3(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n400_), .A2(new_n402_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n455_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n465_), .A3(new_n479_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n482_), .B1(new_n481_), .B2(new_n477_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n455_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n292_), .B(new_n405_), .C1(new_n333_), .C2(new_n328_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(KEYINPUT98), .A3(new_n337_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n342_), .A3(new_n409_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n353_), .B1(new_n279_), .B2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n417_), .B(KEYINPUT27), .C1(new_n497_), .C2(new_n274_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT27), .B1(new_n416_), .B2(new_n417_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n493_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n486_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504_));
  INV_X1    g303(.A(G169gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G197gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G1gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(G8gat), .ZN(new_n512_));
  INV_X1    g311(.A(G8gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(KEYINPUT71), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n510_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n518_), .A3(new_n510_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(G8gat), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n513_), .A2(KEYINPUT71), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n511_), .A2(G8gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(G1gat), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n513_), .A3(new_n519_), .ZN(new_n527_));
  OR2_X1    g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528_));
  INV_X1    g327(.A(G43gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(G43gat), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n531_), .A2(new_n534_), .A3(G50gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(G50gat), .B1(new_n531_), .B2(new_n534_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n521_), .A2(new_n527_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT76), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n521_), .A2(new_n540_), .A3(new_n527_), .A4(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n544_));
  INV_X1    g343(.A(G50gat), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n532_), .A2(new_n533_), .A3(G43gat), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n529_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n531_), .A2(new_n534_), .A3(G50gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(KEYINPUT15), .A3(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n521_), .A2(new_n527_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT77), .ZN(new_n554_));
  AND4_X1   g353(.A1(KEYINPUT78), .A2(new_n542_), .A3(new_n552_), .A4(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT78), .B1(new_n556_), .B2(new_n554_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n521_), .A2(new_n527_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n537_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n542_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(G229gat), .A3(G233gat), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n509_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n542_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(KEYINPUT78), .A3(new_n554_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n563_), .A2(new_n567_), .A3(new_n568_), .A4(new_n509_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n503_), .A2(KEYINPUT100), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT100), .B1(new_n503_), .B2(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n269_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G134gat), .ZN(new_n578_));
  INV_X1    g377(.A(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT36), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n234_), .A2(new_n560_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT68), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT70), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n544_), .A2(new_n550_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n234_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n590_), .A2(KEYINPUT69), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(KEYINPUT69), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n582_), .B(new_n588_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n585_), .A2(new_n586_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n581_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n593_), .A2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n594_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n580_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(KEYINPUT36), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT37), .ZN(new_n604_));
  AND2_X1   g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n243_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n559_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT72), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT16), .B(G183gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT74), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n607_), .A2(KEYINPUT72), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n612_), .B(KEYINPUT17), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n607_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT75), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n604_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT101), .B1(new_n576_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n575_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n268_), .B1(new_n624_), .B2(new_n573_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n626_));
  INV_X1    g425(.A(new_n603_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT37), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n603_), .A2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n621_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(new_n626_), .A3(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n623_), .A2(new_n632_), .A3(new_n510_), .A4(new_n487_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n268_), .B2(new_n571_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n266_), .A2(KEYINPUT103), .A3(new_n572_), .A4(new_n267_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n603_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n620_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n503_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n487_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n633_), .A2(new_n634_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n635_), .A2(new_n643_), .A3(new_n644_), .ZN(G1324gat));
  OAI21_X1  g444(.A(G8gat), .B1(new_n641_), .B2(new_n501_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT39), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n501_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n623_), .A2(new_n632_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n649_), .A3(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  AND2_X1   g453(.A1(new_n623_), .A2(new_n632_), .ZN(new_n655_));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n484_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n639_), .A2(new_n503_), .A3(new_n640_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(new_n484_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(KEYINPUT41), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT41), .B1(new_n661_), .B2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n655_), .A2(new_n666_), .A3(new_n488_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n658_), .B2(new_n488_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(KEYINPUT42), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT42), .B1(new_n670_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n667_), .B1(new_n672_), .B2(new_n673_), .ZN(G1327gat));
  NOR2_X1   g473(.A1(new_n621_), .A2(new_n603_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n269_), .B(new_n675_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n487_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n604_), .B1(new_n486_), .B2(new_n502_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n679_), .B2(KEYINPUT106), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n428_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n428_), .A2(new_n425_), .A3(new_n419_), .A4(new_n418_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n685_), .A2(new_n433_), .A3(new_n417_), .A4(new_n416_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n484_), .B1(new_n686_), .B2(new_n413_), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n687_), .A2(new_n455_), .B1(new_n493_), .B2(new_n501_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n681_), .B(new_n682_), .C1(new_n688_), .C2(new_n604_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n680_), .A2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n620_), .B(KEYINPUT75), .Z(new_n691_));
  AND3_X1   g490(.A1(new_n637_), .A2(new_n638_), .A3(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n690_), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n680_), .A2(new_n689_), .A3(KEYINPUT44), .A4(new_n692_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n642_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n680_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n678_), .B1(new_n697_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n693_), .A2(new_n696_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n501_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n501_), .A2(G36gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT45), .B1(new_n676_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n625_), .A2(new_n711_), .A3(new_n675_), .A4(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n703_), .B1(new_n707_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n501_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n700_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n696_), .B2(new_n693_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT46), .B(new_n713_), .C1(new_n718_), .C2(new_n704_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n719_), .ZN(G1329gat));
  AOI21_X1  g519(.A(new_n529_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n696_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n694_), .A2(new_n695_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n484_), .B(new_n721_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT108), .B(G43gat), .Z(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n676_), .B2(new_n485_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT47), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n729_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n677_), .B2(new_n488_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n455_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n545_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n688_), .A2(new_n572_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n269_), .A2(new_n691_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n642_), .A4(new_n627_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n740_), .A2(KEYINPUT110), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(KEYINPUT110), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n604_), .A3(new_n737_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n743_), .B2(new_n642_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n741_), .A2(new_n742_), .B1(new_n746_), .B2(new_n747_), .ZN(G1332gat));
  OR3_X1    g547(.A1(new_n743_), .A2(G64gat), .A3(new_n501_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n738_), .A2(new_n627_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n716_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G64gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n754_), .A3(G64gat), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n753_), .A2(KEYINPUT48), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT48), .B1(new_n753_), .B2(new_n755_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n749_), .B1(new_n756_), .B2(new_n757_), .ZN(G1333gat));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n484_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G71gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT112), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(G71gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n743_), .A2(G71gat), .A3(new_n485_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n761_), .A2(KEYINPUT49), .A3(new_n763_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(G1334gat));
  OR3_X1    g568(.A1(new_n743_), .A2(G78gat), .A3(new_n455_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n750_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G78gat), .B1(new_n771_), .B2(new_n455_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT50), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT50), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1335gat));
  AND3_X1   g574(.A1(new_n736_), .A2(new_n268_), .A3(new_n675_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n487_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n572_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n691_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n691_), .B2(new_n778_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n690_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n487_), .A2(G85gat), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT114), .Z(new_n785_));
  AOI21_X1  g584(.A(new_n777_), .B1(new_n783_), .B2(new_n785_), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n690_), .A2(new_n716_), .A3(new_n782_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G92gat), .ZN(new_n788_));
  INV_X1    g587(.A(G92gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n776_), .A2(new_n789_), .A3(new_n716_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT115), .ZN(G1337gat));
  NAND3_X1  g591(.A1(new_n690_), .A2(new_n484_), .A3(new_n782_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(G99gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n776_), .A2(new_n229_), .A3(new_n484_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g596(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n680_), .A2(new_n782_), .A3(new_n689_), .A4(new_n488_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G106gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT52), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n776_), .A2(new_n209_), .A3(new_n488_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n800_), .A2(KEYINPUT52), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n799_), .B2(G106gat), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n798_), .B(new_n802_), .C1(new_n804_), .C2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n803_), .A2(new_n808_), .ZN(G1339gat));
  NOR2_X1   g608(.A1(new_n716_), .A2(new_n642_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n492_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(new_n250_), .B2(new_n251_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n817_), .B(new_n254_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n247_), .A2(new_n254_), .A3(new_n249_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n816_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n821_), .B2(new_n261_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n252_), .A2(new_n817_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n250_), .A2(KEYINPUT55), .A3(new_n251_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n819_), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n262_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n264_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n563_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n508_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n830_), .B2(new_n569_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n562_), .A2(new_n554_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n556_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n832_), .B(new_n508_), .C1(new_n833_), .C2(new_n554_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n569_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n569_), .A2(new_n837_), .A3(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n263_), .A2(new_n264_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n827_), .A2(new_n831_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n814_), .B(KEYINPUT57), .C1(new_n841_), .C2(new_n627_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n821_), .A2(new_n815_), .A3(new_n261_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n262_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n831_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n838_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n837_), .B1(new_n569_), .B2(new_n834_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n840_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n627_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n843_), .B1(new_n850_), .B2(KEYINPUT118), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n842_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n828_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT58), .B1(new_n853_), .B2(new_n839_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n604_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n839_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n640_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n266_), .A2(new_n571_), .A3(new_n267_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n631_), .B2(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n622_), .A2(KEYINPUT54), .A3(new_n861_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n572_), .B(new_n813_), .C1(new_n859_), .C2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n375_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n870_));
  AOI21_X1  g669(.A(new_n621_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n813_), .B(new_n870_), .C1(new_n871_), .C2(new_n865_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n571_), .A2(new_n375_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n264_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n265_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n603_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n877_), .B2(new_n814_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n850_), .A2(KEYINPUT118), .A3(new_n843_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n858_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n620_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n631_), .A2(new_n860_), .A3(new_n862_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n622_), .B2(new_n861_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n812_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n872_), .B(new_n873_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n866_), .A2(KEYINPUT119), .A3(new_n375_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n869_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT121), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n869_), .A2(new_n887_), .A3(new_n891_), .A4(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1340gat));
  OAI21_X1  g692(.A(new_n872_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G120gat), .B1(new_n894_), .B2(new_n269_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n381_), .B1(new_n269_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n885_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n381_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1341gat));
  AOI21_X1  g697(.A(G127gat), .B1(new_n885_), .B2(new_n621_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n894_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT122), .B(G127gat), .Z(new_n901_));
  NOR2_X1   g700(.A1(new_n620_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(G1342gat));
  AOI21_X1  g702(.A(G134gat), .B1(new_n885_), .B2(new_n627_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n604_), .A2(new_n376_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n900_), .B2(new_n905_), .ZN(G1343gat));
  NOR2_X1   g705(.A1(new_n859_), .A2(new_n865_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n489_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n810_), .A2(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT123), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n572_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n268_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g714(.A1(new_n907_), .A2(new_n691_), .A3(new_n910_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n911_), .A2(G162gat), .A3(new_n856_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n911_), .A2(new_n627_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n579_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n921_), .A2(KEYINPUT124), .A3(new_n579_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n920_), .B1(new_n924_), .B2(new_n925_), .ZN(G1347gat));
  AND3_X1   g725(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n839_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n854_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n851_), .A2(new_n842_), .B1(new_n928_), .B2(new_n856_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n884_), .B1(new_n929_), .B2(new_n621_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n501_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n505_), .B1(new_n932_), .B2(new_n572_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n933_), .A2(KEYINPUT62), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n572_), .A3(new_n321_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(KEYINPUT62), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n936_), .ZN(G1348gat));
  OAI21_X1  g736(.A(new_n884_), .B1(new_n929_), .B2(new_n640_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n501_), .A2(new_n487_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n938_), .A2(new_n455_), .A3(new_n484_), .A4(new_n939_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n940_), .A2(new_n322_), .A3(new_n269_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G176gat), .B1(new_n932_), .B2(new_n268_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1349gat));
  OAI211_X1 g742(.A(new_n621_), .B(new_n931_), .C1(new_n859_), .C2(new_n865_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n938_), .A2(KEYINPUT125), .A3(new_n621_), .A4(new_n931_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n946_), .A2(new_n317_), .A3(new_n947_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n932_), .A2(new_n332_), .A3(new_n330_), .A4(new_n640_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT126), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n948_), .A2(new_n949_), .A3(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n932_), .A2(new_n627_), .A3(new_n347_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n932_), .A2(new_n856_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n955_), .B1(new_n957_), .B2(new_n318_), .ZN(G1351gat));
  NAND4_X1  g757(.A1(new_n938_), .A2(new_n572_), .A3(new_n908_), .A4(new_n939_), .ZN(new_n959_));
  OR3_X1    g758(.A1(new_n959_), .A2(KEYINPUT127), .A3(new_n507_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n507_), .ZN(new_n961_));
  OAI21_X1  g760(.A(KEYINPUT127), .B1(new_n959_), .B2(new_n507_), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n960_), .A2(new_n961_), .A3(new_n962_), .ZN(G1352gat));
  NAND3_X1  g762(.A1(new_n938_), .A2(new_n908_), .A3(new_n939_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n269_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(new_n286_), .ZN(G1353gat));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AND2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  NOR4_X1   g767(.A1(new_n964_), .A2(new_n620_), .A3(new_n967_), .A4(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n964_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n640_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n969_), .B1(new_n971_), .B2(new_n967_), .ZN(G1354gat));
  AOI21_X1  g771(.A(G218gat), .B1(new_n970_), .B2(new_n627_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n964_), .A2(new_n604_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(G218gat), .B2(new_n974_), .ZN(G1355gat));
endmodule


