//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_, new_n967_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT2), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G141gat), .A3(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OAI22_X1  g006(.A1(KEYINPUT85), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G155gat), .ZN(new_n214_));
  INV_X1    g013(.A(G162gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT83), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT84), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT84), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G155gat), .A3(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n219_), .A2(new_n224_), .A3(KEYINPUT86), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT86), .B1(new_n219_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n213_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n210_), .A2(new_n211_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(new_n223_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n219_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n203_), .B(new_n228_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G134gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G127gat), .ZN(new_n235_));
  INV_X1    g034(.A(G127gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G134gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT82), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT82), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT82), .B1(new_n235_), .B2(new_n237_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n227_), .A2(new_n233_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n202_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n243_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n207_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n219_), .A2(new_n224_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n219_), .A2(new_n224_), .A3(KEYINPUT86), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n252_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n228_), .A2(new_n203_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n230_), .A2(new_n219_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n232_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n251_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n247_), .A2(new_n243_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(new_n227_), .A3(new_n233_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(KEYINPUT4), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n250_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n202_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT0), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G57gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G85gat), .ZN(new_n272_));
  INV_X1    g071(.A(G57gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n270_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G85gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n266_), .A2(new_n267_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G15gat), .B(G43gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT81), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT24), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G190gat), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n293_), .A2(KEYINPUT78), .A3(KEYINPUT26), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT26), .B1(new_n293_), .B2(KEYINPUT78), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G183gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT25), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G183gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT77), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(KEYINPUT77), .B2(new_n298_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n292_), .B1(new_n296_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT79), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT79), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n305_), .A2(new_n307_), .A3(KEYINPUT23), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n297_), .A2(new_n293_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G169gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT22), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G169gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n289_), .B1(new_n321_), .B2(G176gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n303_), .A2(new_n311_), .B1(new_n316_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n290_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n291_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n287_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n299_), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT25), .B(G183gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(KEYINPUT77), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n294_), .A2(new_n295_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n330_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n309_), .A2(new_n310_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n312_), .A2(new_n313_), .B1(new_n297_), .B2(new_n293_), .ZN(new_n337_));
  OAI22_X1  g136(.A1(new_n335_), .A2(new_n336_), .B1(new_n337_), .B2(new_n322_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(new_n325_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n286_), .B1(new_n327_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n286_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n324_), .A2(new_n326_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n325_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n251_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n340_), .A2(new_n344_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT31), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n263_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT29), .B1(new_n257_), .B2(new_n261_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT89), .ZN(new_n355_));
  INV_X1    g154(.A(G211gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(G218gat), .ZN(new_n357_));
  INV_X1    g156(.A(G218gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(G211gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n355_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(G211gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(G218gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT89), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G197gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT87), .B1(new_n365_), .B2(G204gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367_));
  INV_X1    g166(.A(G204gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(G197gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(G204gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n366_), .A2(new_n369_), .A3(KEYINPUT90), .A4(new_n370_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n364_), .A2(new_n373_), .A3(KEYINPUT21), .A4(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n370_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n365_), .A2(G204gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT21), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n357_), .A2(new_n359_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n380_));
  OAI211_X1 g179(.A(new_n378_), .B(new_n379_), .C1(new_n371_), .C2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n354_), .B(new_n382_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n383_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n384_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n375_), .A2(new_n381_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n386_), .B(new_n387_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n385_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT92), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(new_n391_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n392_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n385_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n227_), .A2(new_n233_), .A3(new_n388_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT28), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n227_), .A2(new_n404_), .A3(new_n388_), .A4(new_n233_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G22gat), .B(G50gat), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n396_), .A2(new_n401_), .A3(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n410_), .B(KEYINPUT92), .C1(new_n394_), .C2(new_n395_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n353_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT97), .ZN(new_n415_));
  AND2_X1   g214(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n289_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT95), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n289_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n329_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n293_), .A2(KEYINPUT26), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT26), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G190gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT93), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n332_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n416_), .A2(new_n417_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n312_), .A2(new_n313_), .B1(new_n430_), .B2(new_n291_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n319_), .A2(G169gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n317_), .A2(KEYINPUT22), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT96), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G176gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n318_), .A2(new_n320_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n309_), .A2(new_n315_), .A3(new_n310_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n289_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n390_), .A2(new_n415_), .A3(new_n432_), .A4(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n432_), .A2(new_n381_), .A3(new_n375_), .A4(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT97), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT19), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n338_), .B2(new_n382_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n442_), .A2(new_n444_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n311_), .B(new_n330_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n316_), .A2(new_n323_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n381_), .A4(new_n375_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT20), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n432_), .A2(new_n441_), .B1(new_n375_), .B2(new_n381_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n446_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G8gat), .B(G36gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT18), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n450_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT101), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n450_), .A2(new_n461_), .A3(new_n456_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n461_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT101), .B(new_n466_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n464_), .A2(KEYINPUT27), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT100), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n432_), .A2(new_n441_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n382_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n476_), .A2(KEYINPUT20), .A3(new_n453_), .A4(new_n447_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT98), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n448_), .B1(new_n390_), .B2(new_n324_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT98), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n447_), .A4(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n449_), .A2(new_n443_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n478_), .A2(new_n481_), .B1(new_n446_), .B2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n473_), .B(new_n474_), .C1(new_n461_), .C2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n446_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n461_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n464_), .A2(KEYINPUT27), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT100), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  AND4_X1   g289(.A1(new_n280_), .A2(new_n414_), .A3(new_n472_), .A4(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n412_), .A2(new_n413_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n472_), .A2(new_n490_), .A3(new_n492_), .A4(new_n280_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n262_), .A2(KEYINPUT4), .A3(new_n264_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n202_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n262_), .B2(KEYINPUT4), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n267_), .B(new_n277_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT33), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n266_), .A2(KEYINPUT33), .A3(new_n267_), .A4(new_n277_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n277_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n262_), .A2(new_n264_), .A3(new_n495_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n202_), .B1(new_n262_), .B2(KEYINPUT4), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n501_), .B(new_n502_), .C1(new_n494_), .C2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n461_), .A2(KEYINPUT32), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n450_), .A2(new_n456_), .A3(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n509_));
  OAI22_X1  g308(.A1(new_n465_), .A2(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n412_), .A2(new_n413_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT99), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT99), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n493_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n491_), .B1(new_n516_), .B2(new_n353_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G1gat), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G29gat), .B(G36gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n524_), .A2(new_n531_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n531_), .B(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n535_), .B2(new_n524_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  MUX2_X1   g336(.A(new_n532_), .B(new_n536_), .S(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(KEYINPUT76), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT74), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT75), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G169gat), .B(G197gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n540_), .A2(new_n545_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(G92gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n275_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(G99gat), .A3(G106gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n558_));
  NAND2_X1  g357(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n559_));
  INV_X1    g358(.A(G99gat), .ZN(new_n560_));
  INV_X1    g359(.A(G106gat), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n558_), .B(new_n559_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  OR3_X1    g362(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n555_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT8), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n555_), .A2(KEYINPUT8), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n557_), .B(new_n562_), .C1(KEYINPUT65), .C2(new_n566_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n566_), .A2(KEYINPUT65), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n553_), .A2(KEYINPUT9), .A3(new_n554_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n554_), .A2(KEYINPUT9), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT10), .B(G99gat), .Z(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n561_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n563_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n569_), .A2(new_n573_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT11), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584_));
  INV_X1    g383(.A(KEYINPUT66), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT66), .ZN(new_n588_));
  AOI211_X1 g387(.A(new_n582_), .B(new_n583_), .C1(new_n586_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n583_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n588_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(KEYINPUT11), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n586_), .A2(new_n582_), .A3(new_n588_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n581_), .A2(KEYINPUT67), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT67), .B1(new_n581_), .B2(new_n594_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n581_), .A2(new_n594_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n551_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n550_), .B1(new_n581_), .B2(new_n594_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT69), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n594_), .A2(KEYINPUT12), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT68), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n581_), .A2(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n567_), .A2(new_n568_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(KEYINPUT68), .A3(new_n573_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT12), .B1(new_n581_), .B2(new_n594_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT69), .B(new_n550_), .C1(new_n581_), .C2(new_n594_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n602_), .A2(new_n608_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT70), .ZN(new_n615_));
  XOR2_X1   g414(.A(G176gat), .B(G204gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n599_), .A2(new_n612_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT72), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT72), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n599_), .A2(new_n612_), .A3(new_n620_), .A4(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n599_), .A2(new_n612_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n617_), .B(KEYINPUT71), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n622_), .A2(KEYINPUT13), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT13), .B1(new_n622_), .B2(new_n625_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n517_), .A2(new_n549_), .A3(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n581_), .A2(new_n604_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT68), .B1(new_n606_), .B2(new_n573_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n535_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n581_), .A2(new_n531_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT35), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n634_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n633_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n635_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643_));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(KEYINPUT36), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n633_), .B(new_n639_), .C1(new_n635_), .C2(new_n638_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n642_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n645_), .B(KEYINPUT36), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n642_), .B2(new_n648_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT37), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n524_), .B(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(new_n594_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G127gat), .B(G155gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT16), .ZN(new_n662_));
  XOR2_X1   g461(.A(G183gat), .B(G211gat), .Z(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT17), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n664_), .A2(new_n665_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n660_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n666_), .B2(new_n660_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n657_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n629_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n280_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n629_), .A2(KEYINPUT102), .A3(new_n671_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n674_), .A2(new_n519_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n677_), .A2(KEYINPUT103), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(KEYINPUT103), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(KEYINPUT38), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT104), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT38), .B1(new_n678_), .B2(new_n679_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n517_), .A2(new_n653_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n628_), .A2(new_n549_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n669_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n519_), .B1(new_n686_), .B2(new_n675_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n682_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n688_), .ZN(G1324gat));
  INV_X1    g488(.A(new_n472_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n490_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n520_), .B1(new_n686_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT105), .B1(new_n695_), .B2(KEYINPUT39), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT39), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n696_), .B(new_n699_), .C1(new_n698_), .C2(new_n694_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n674_), .A2(new_n676_), .A3(new_n520_), .A4(new_n693_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT40), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1325gat));
  INV_X1    g505(.A(G15gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n353_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n686_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n707_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n711_), .B(new_n712_), .C1(new_n672_), .C2(new_n713_), .ZN(G1326gat));
  INV_X1    g513(.A(G22gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n686_), .B2(new_n492_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT42), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n672_), .A2(G22gat), .A3(new_n511_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1327gat));
  INV_X1    g518(.A(new_n653_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n669_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n629_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G29gat), .B1(new_n723_), .B2(new_n675_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n657_), .ZN(new_n725_));
  NOR4_X1   g524(.A1(new_n517_), .A2(new_n725_), .A3(KEYINPUT106), .A4(KEYINPUT43), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n517_), .B2(new_n725_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n517_), .A2(KEYINPUT43), .A3(new_n725_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n684_), .A2(new_n670_), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n734_), .A2(G29gat), .A3(new_n675_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n724_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  XOR2_X1   g536(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n692_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(G36gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n739_), .B1(new_n723_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n745_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n722_), .A3(new_n738_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n746_), .A2(new_n748_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n734_), .A2(new_n693_), .A3(new_n736_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G36gat), .ZN(new_n751_));
  AND2_X1   g550(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1329gat));
  NAND3_X1  g552(.A1(new_n734_), .A2(G43gat), .A3(new_n708_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n736_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n722_), .A2(new_n353_), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n754_), .A2(new_n755_), .B1(G43gat), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g557(.A(G50gat), .B1(new_n723_), .B2(new_n492_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n734_), .A2(G50gat), .A3(new_n492_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n736_), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n626_), .A2(new_n627_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n517_), .A2(new_n548_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n671_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n273_), .A3(new_n675_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n628_), .A2(new_n669_), .A3(new_n549_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n683_), .A2(new_n280_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n768_), .B2(new_n273_), .ZN(G1332gat));
  INV_X1    g568(.A(G64gat), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n683_), .A2(new_n767_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n743_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT48), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n743_), .A2(new_n770_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT110), .Z(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n764_), .B2(new_n775_), .ZN(G1333gat));
  INV_X1    g575(.A(G71gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n771_), .B2(new_n708_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT49), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n777_), .A3(new_n708_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1334gat));
  INV_X1    g580(.A(G78gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n771_), .B2(new_n492_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT50), .Z(new_n784_));
  NAND3_X1  g583(.A1(new_n765_), .A2(new_n782_), .A3(new_n492_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1335gat));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n628_), .A2(new_n670_), .A3(new_n549_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n731_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n788_), .B(KEYINPUT112), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n517_), .A2(KEYINPUT43), .A3(new_n725_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n728_), .B2(new_n727_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT113), .B(new_n792_), .C1(new_n794_), .C2(new_n726_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n280_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n763_), .A2(new_n721_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT111), .Z(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n275_), .A3(new_n675_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n796_), .B2(new_n744_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n552_), .A3(new_n693_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1337gat));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n577_), .A3(new_n708_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n353_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n560_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n492_), .B(new_n792_), .C1(new_n794_), .C2(new_n726_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(G106gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n810_), .B2(G106gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n731_), .A2(new_n511_), .A3(new_n790_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT114), .B1(new_n815_), .B2(new_n561_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n810_), .A2(new_n811_), .A3(G106gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(KEYINPUT52), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n799_), .A2(new_n561_), .A3(new_n492_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT53), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n814_), .A2(new_n818_), .A3(new_n819_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1339gat));
  NAND2_X1  g623(.A1(new_n622_), .A2(new_n548_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT116), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n602_), .A2(new_n611_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n609_), .B1(new_n632_), .B2(new_n603_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(KEYINPUT55), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n612_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n608_), .A2(new_n610_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n551_), .B1(new_n832_), .B2(new_n598_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n624_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n624_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n622_), .A2(new_n548_), .A3(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n826_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n622_), .A2(new_n625_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n538_), .A2(new_n545_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n536_), .A2(G229gat), .A3(G233gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n532_), .A2(new_n537_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n545_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n653_), .B1(new_n842_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n622_), .A2(new_n849_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT117), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n848_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n853_), .A2(new_n839_), .A3(KEYINPUT58), .A4(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n657_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n837_), .A2(new_n838_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT58), .B1(new_n859_), .B2(new_n853_), .ZN(new_n860_));
  OAI22_X1  g659(.A1(new_n851_), .A2(KEYINPUT57), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n862_), .B(new_n653_), .C1(new_n842_), .C2(new_n850_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n670_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  AND4_X1   g663(.A1(new_n669_), .A2(new_n654_), .A3(new_n656_), .A4(new_n549_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n762_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT115), .B1(new_n866_), .B2(KEYINPUT54), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n865_), .A2(new_n762_), .A3(new_n868_), .A4(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n866_), .A2(KEYINPUT54), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n692_), .A2(new_n708_), .A3(new_n675_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n511_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT59), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n873_), .A2(new_n511_), .A3(new_n875_), .A4(new_n879_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n548_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G113gat), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n876_), .A2(G113gat), .A3(new_n549_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1340gat));
  NAND3_X1  g684(.A1(new_n877_), .A2(new_n628_), .A3(new_n880_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT119), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G120gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(KEYINPUT119), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n762_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n891_));
  OAI22_X1  g690(.A1(new_n888_), .A2(new_n889_), .B1(new_n876_), .B2(new_n891_), .ZN(G1341gat));
  OAI21_X1  g691(.A(new_n236_), .B1(new_n876_), .B2(new_n670_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT120), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n670_), .A2(new_n236_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n881_), .B2(new_n895_), .ZN(G1342gat));
  AOI211_X1 g695(.A(new_n492_), .B(new_n874_), .C1(new_n864_), .C2(new_n872_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n880_), .B(new_n657_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G134gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(new_n234_), .A3(new_n653_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(KEYINPUT121), .A3(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1343gat));
  AOI211_X1 g705(.A(new_n708_), .B(new_n511_), .C1(new_n864_), .C2(new_n872_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n743_), .A2(new_n280_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n549_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n210_), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n762_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n211_), .ZN(G1345gat));
  NOR2_X1   g712(.A1(new_n909_), .A2(new_n670_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT61), .B(G155gat), .Z(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  OAI21_X1  g715(.A(new_n215_), .B1(new_n909_), .B2(new_n720_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n657_), .A2(G162gat), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT122), .Z(new_n919_));
  NAND3_X1  g718(.A1(new_n907_), .A2(new_n908_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n917_), .A2(KEYINPUT123), .A3(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1347gat));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n492_), .B1(new_n864_), .B2(new_n872_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n744_), .A2(new_n675_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n708_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n549_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n926_), .B1(new_n932_), .B2(new_n317_), .ZN(new_n933_));
  OAI211_X1 g732(.A(KEYINPUT62), .B(G169gat), .C1(new_n931_), .C2(new_n549_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(G1348gat));
  NAND2_X1  g735(.A1(new_n873_), .A2(new_n511_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(KEYINPUT124), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n927_), .A2(new_n939_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n929_), .A2(new_n436_), .A3(new_n762_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n436_), .B1(new_n931_), .B2(new_n762_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1349gat));
  NOR3_X1   g745(.A1(new_n931_), .A2(new_n670_), .A3(new_n332_), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n938_), .A2(new_n669_), .A3(new_n930_), .A4(new_n940_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n297_), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n931_), .B2(new_n725_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n653_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n931_), .B2(new_n951_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT126), .ZN(G1351gat));
  NAND2_X1  g752(.A1(new_n907_), .A2(new_n928_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n549_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(new_n365_), .ZN(G1352gat));
  NOR2_X1   g755(.A1(new_n954_), .A2(new_n762_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(new_n368_), .ZN(G1353gat));
  NOR2_X1   g757(.A1(new_n954_), .A2(new_n670_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  AND2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n959_), .B1(new_n960_), .B2(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n962_), .B1(new_n959_), .B2(new_n960_), .ZN(G1354gat));
  NOR3_X1   g762(.A1(new_n954_), .A2(new_n358_), .A3(new_n725_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n954_), .A2(new_n720_), .ZN(new_n965_));
  OR2_X1    g764(.A1(new_n965_), .A2(KEYINPUT127), .ZN(new_n966_));
  AOI21_X1  g765(.A(G218gat), .B1(new_n965_), .B2(KEYINPUT127), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n964_), .B1(new_n966_), .B2(new_n967_), .ZN(G1355gat));
endmodule


