//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT82), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT3), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n223_), .A2(new_n213_), .A3(new_n214_), .A4(KEYINPUT82), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n204_), .A2(new_n203_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT83), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(new_n229_), .A3(new_n226_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n217_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n202_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G211gat), .B(G218gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G197gat), .B(G204gat), .Z(new_n235_));
  AOI21_X1  g034(.A(new_n234_), .B1(KEYINPUT21), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G204gat), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n237_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT86), .B1(new_n237_), .B2(G197gat), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n238_), .A2(new_n239_), .B1(G197gat), .B2(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n236_), .B1(KEYINPUT21), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT89), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(KEYINPUT21), .A3(new_n234_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n225_), .A2(new_n229_), .A3(new_n226_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n229_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n233_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n241_), .A2(new_n243_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(new_n256_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n250_), .B2(KEYINPUT29), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(KEYINPUT87), .A3(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G78gat), .B(G106gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT90), .Z(new_n264_));
  AND3_X1   g063(.A1(new_n255_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n255_), .B2(new_n262_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT92), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n255_), .A2(new_n262_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n264_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n255_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G22gat), .B(G50gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n231_), .A2(new_n232_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT84), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(KEYINPUT84), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n277_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n278_), .A2(KEYINPUT84), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT91), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(new_n272_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n267_), .A2(new_n273_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n287_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT92), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n271_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(G127gat), .A2(G134gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT78), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(G127gat), .A2(G134gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G127gat), .A2(G134gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT78), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G120gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n296_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n247_), .B(new_n303_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n228_), .A2(new_n230_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n307_), .A2(KEYINPUT98), .A3(new_n247_), .A4(new_n303_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(new_n299_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n300_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n296_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT79), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n250_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT97), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n250_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n309_), .A2(KEYINPUT4), .A3(new_n319_), .A4(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n318_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n309_), .A2(new_n323_), .A3(new_n319_), .A4(new_n321_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT0), .B(G57gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G85gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(G1gat), .B(G29gat), .Z(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT33), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n334_), .A2(KEYINPUT99), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n334_), .B2(KEYINPUT99), .ZN(new_n337_));
  INV_X1    g136(.A(new_n323_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n322_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n309_), .A2(new_n338_), .A3(new_n319_), .A4(new_n321_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n332_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT18), .B(G64gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT23), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  INV_X1    g148(.A(G176gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n351_), .A2(KEYINPUT24), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT25), .B(G183gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(KEYINPUT24), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT76), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(KEYINPUT76), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n353_), .A2(new_n356_), .A3(new_n359_), .A4(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n348_), .B1(G183gat), .B2(G190gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT22), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(KEYINPUT77), .B2(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n350_), .B1(new_n365_), .B2(KEYINPUT22), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n362_), .B(new_n357_), .C1(new_n364_), .C2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n361_), .A2(new_n367_), .A3(new_n241_), .A4(new_n243_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT96), .ZN(new_n369_));
  INV_X1    g168(.A(new_n357_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(G169gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n349_), .A2(KEYINPUT22), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n350_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT95), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n357_), .A2(KEYINPUT95), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n369_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G169gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT95), .B1(new_n379_), .B2(new_n350_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT96), .B(new_n378_), .C1(new_n380_), .C2(new_n370_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n353_), .A2(new_n383_), .A3(new_n356_), .A4(new_n358_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n356_), .A2(new_n348_), .A3(new_n352_), .A4(new_n358_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT94), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n382_), .A2(new_n362_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n256_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT20), .B(new_n368_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(KEYINPUT93), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n388_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n391_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n361_), .A2(new_n367_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n397_), .B2(new_n256_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n346_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(new_n346_), .A3(new_n399_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n342_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n336_), .A2(new_n337_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n393_), .A2(new_n399_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n389_), .A2(new_n392_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n382_), .A2(new_n362_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n385_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n395_), .B1(new_n410_), .B2(new_n398_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n406_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n334_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n333_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n407_), .B(new_n412_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n288_), .B(new_n292_), .C1(new_n404_), .C2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n413_), .A2(new_n414_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT27), .ZN(new_n419_));
  INV_X1    g218(.A(new_n402_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(new_n400_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n408_), .A2(new_n411_), .ZN(new_n422_));
  OAI211_X1 g221(.A(KEYINPUT27), .B(new_n402_), .C1(new_n422_), .C2(new_n346_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n267_), .A2(new_n273_), .A3(new_n287_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n287_), .B1(new_n267_), .B2(new_n273_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n418_), .B(new_n424_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n417_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n311_), .A2(new_n316_), .A3(new_n433_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n361_), .A3(new_n367_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n397_), .B1(new_n438_), .B2(new_n434_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT31), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n432_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n439_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n441_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n431_), .A3(new_n443_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT80), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n425_), .A2(new_n426_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n414_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n450_), .A2(new_n454_), .A3(new_n334_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n453_), .A2(KEYINPUT100), .A3(new_n424_), .A4(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n292_), .A2(new_n288_), .A3(new_n424_), .A4(new_n455_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n428_), .A2(new_n452_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G57gat), .B(G64gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT64), .ZN(new_n462_));
  INV_X1    g261(.A(G57gat), .ZN(new_n463_));
  INV_X1    g262(.A(G64gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G57gat), .A2(G64gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n462_), .A2(new_n473_), .A3(new_n468_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(KEYINPUT11), .A3(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT10), .B(G99gat), .Z(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G85gat), .B(G92gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT9), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G85gat), .A3(G92gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n480_), .A2(new_n482_), .A3(new_n484_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n479_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n493_), .A2(new_n487_), .A3(new_n488_), .A4(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n481_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(KEYINPUT8), .A3(new_n481_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n477_), .A2(new_n490_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n490_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(KEYINPUT12), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(KEYINPUT12), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n503_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G120gat), .B(G148gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(new_n237_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT5), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(new_n350_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n512_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n508_), .B(new_n511_), .C1(KEYINPUT65), .C2(new_n517_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT13), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n349_), .ZN(new_n524_));
  INV_X1    g323(.A(G197gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527_));
  INV_X1    g326(.A(G1gat), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G8gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G29gat), .B(G36gat), .Z(new_n534_));
  INV_X1    g333(.A(G43gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G29gat), .B(G36gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G43gat), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(G50gat), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(G50gat), .B1(new_n536_), .B2(new_n538_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n538_), .ZN(new_n543_));
  INV_X1    g342(.A(G50gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(G50gat), .A3(new_n538_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT15), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n533_), .B1(new_n542_), .B2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n531_), .B(new_n532_), .Z(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n546_), .A3(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT74), .Z(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n533_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n550_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n551_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n545_), .A2(new_n546_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(KEYINPUT73), .A3(new_n533_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n557_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n526_), .B1(new_n554_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n526_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n553_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(KEYINPUT75), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n567_), .B(new_n526_), .C1(new_n554_), .C2(new_n561_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n522_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n460_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n502_), .B1(new_n542_), .B2(new_n547_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT66), .B(KEYINPUT34), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT67), .ZN(new_n575_));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n559_), .A2(new_n502_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n573_), .A2(KEYINPUT35), .A3(new_n580_), .A4(new_n582_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G134gat), .ZN(new_n587_));
  INV_X1    g386(.A(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(new_n590_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n584_), .B(new_n585_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n592_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n572_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT70), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(KEYINPUT68), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n584_), .A2(new_n585_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n591_), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT69), .B1(new_n601_), .B2(new_n594_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT68), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT70), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n594_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n603_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n599_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n599_), .B2(new_n604_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(G231gat), .ZN(new_n611_));
  INV_X1    g410(.A(G233gat), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n477_), .A2(new_n549_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n477_), .A2(new_n549_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n613_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n613_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n614_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n621_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n617_), .B(new_n620_), .C1(new_n627_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT72), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT72), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n630_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n610_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n571_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n418_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n528_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n635_), .A2(new_n606_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n571_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n418_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1324gat));
  OAI21_X1  g443(.A(KEYINPUT101), .B1(new_n642_), .B2(new_n424_), .ZN(new_n645_));
  NOR4_X1   g444(.A1(new_n460_), .A2(new_n635_), .A3(new_n606_), .A4(new_n570_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(new_n424_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(G8gat), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT39), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n637_), .A2(new_n529_), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(KEYINPUT40), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n646_), .B2(new_n451_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n637_), .A2(new_n658_), .A3(new_n451_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1326gat));
  OAI21_X1  g461(.A(G22gat), .B1(new_n642_), .B2(new_n453_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT102), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n665_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n453_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n637_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n666_), .B(new_n667_), .C1(G22gat), .C2(new_n669_), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n599_), .A2(new_n604_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n607_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n599_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n456_), .A2(new_n459_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n451_), .B1(new_n417_), .B2(new_n427_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n677_), .B(new_n610_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n522_), .A2(new_n635_), .A3(new_n569_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT104), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n428_), .A2(new_n452_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n456_), .A2(new_n459_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n677_), .B1(new_n692_), .B2(new_n610_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT43), .B(new_n675_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n683_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(KEYINPUT103), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n689_), .A2(new_n700_), .A3(new_n638_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G29gat), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n635_), .A2(new_n606_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT105), .Z(new_n704_));
  NAND2_X1  g503(.A1(new_n571_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n418_), .A2(G29gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT106), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n705_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT103), .B1(new_n695_), .B2(new_n696_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n686_), .A2(new_n698_), .A3(KEYINPUT44), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n648_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n688_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n687_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G36gat), .B1(new_n715_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n705_), .A2(G36gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n648_), .ZN(new_n723_));
  NOR4_X1   g522(.A1(new_n705_), .A2(G36gat), .A3(new_n424_), .A4(new_n720_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n723_), .A2(new_n724_), .B1(KEYINPUT108), .B2(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n712_), .B1(new_n719_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G36gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n424_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n689_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n730_), .A2(new_n711_), .A3(new_n725_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1329gat));
  OAI21_X1  g531(.A(new_n535_), .B1(new_n705_), .B2(new_n452_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n689_), .A2(G43gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n700_), .A2(new_n450_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n733_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1330gat));
  NAND3_X1  g539(.A1(new_n689_), .A2(new_n700_), .A3(new_n668_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G50gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n453_), .A2(G50gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT110), .ZN(new_n746_));
  OAI22_X1  g545(.A1(new_n743_), .A2(new_n744_), .B1(new_n705_), .B2(new_n746_), .ZN(G1331gat));
  INV_X1    g546(.A(KEYINPUT13), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n521_), .B(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n636_), .A2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT111), .Z(new_n751_));
  NAND2_X1  g550(.A1(new_n566_), .A2(new_n568_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n692_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT112), .ZN(new_n754_));
  AOI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n638_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n460_), .A2(new_n569_), .A3(new_n522_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n641_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n638_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(G57gat), .B2(new_n758_), .ZN(G1332gat));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n464_), .A3(new_n648_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n464_), .B1(new_n757_), .B2(new_n648_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT48), .Z(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n764_), .A3(new_n451_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n757_), .B2(new_n451_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT49), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1334gat));
  INV_X1    g567(.A(G78gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n754_), .A2(new_n769_), .A3(new_n668_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n757_), .B2(new_n668_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT50), .Z(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n756_), .A2(new_n704_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(G85gat), .A3(new_n418_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n522_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n635_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n569_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n638_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n775_), .B1(new_n780_), .B2(G85gat), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT113), .ZN(G1336gat));
  INV_X1    g581(.A(new_n774_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G92gat), .B1(new_n783_), .B2(new_n648_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n648_), .A2(G92gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT114), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n779_), .B2(new_n786_), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n776_), .A2(new_n451_), .A3(new_n778_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G99gat), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT51), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n450_), .A2(new_n478_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n789_), .B(new_n791_), .C1(new_n774_), .C2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n790_), .A2(KEYINPUT51), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n793_), .B(new_n794_), .Z(G1338gat));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n479_), .A3(new_n668_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n776_), .A2(new_n668_), .A3(new_n778_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1339gat));
  INV_X1    g602(.A(G113gat), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT55), .B(new_n510_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n806_), .A2(new_n807_), .B1(new_n507_), .B2(new_n506_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n518_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n557_), .A2(new_n560_), .A3(new_n552_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n548_), .A2(new_n550_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n811_), .B(new_n526_), .C1(new_n812_), .C2(new_n552_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n565_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n512_), .A2(new_n518_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n808_), .A2(new_n818_), .A3(new_n518_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n810_), .A2(new_n815_), .A3(new_n817_), .A4(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n816_), .B1(new_n809_), .B2(KEYINPUT56), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n815_), .A4(new_n819_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n822_), .A2(new_n673_), .A3(new_n674_), .A4(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n814_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n808_), .A2(new_n518_), .A3(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(new_n569_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n828_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n816_), .B1(new_n809_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n827_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n826_), .B1(new_n833_), .B2(new_n606_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n809_), .A2(new_n831_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(new_n569_), .A3(new_n829_), .A4(new_n817_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n827_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n606_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n825_), .A2(new_n834_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n635_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n749_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n635_), .B2(new_n569_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n632_), .A2(new_n752_), .A3(KEYINPUT117), .A4(new_n634_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n845_), .A2(new_n846_), .A3(KEYINPUT54), .A4(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n850_), .B(new_n522_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n846_), .A2(KEYINPUT54), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n846_), .A2(KEYINPUT54), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n841_), .A2(KEYINPUT122), .A3(new_n635_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n844_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n453_), .A2(new_n638_), .A3(new_n424_), .A4(new_n450_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n862_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n859_), .A2(new_n860_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n825_), .A2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n610_), .A2(KEYINPUT120), .A3(new_n822_), .A4(new_n824_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n840_), .A4(new_n834_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n856_), .B1(new_n871_), .B2(new_n635_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT59), .B1(new_n872_), .B2(new_n865_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n867_), .A2(KEYINPUT123), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n859_), .A2(new_n866_), .A3(new_n875_), .A4(new_n860_), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n804_), .B(new_n752_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n872_), .A2(new_n865_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G113gat), .B1(new_n878_), .B2(new_n569_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n874_), .A2(new_n876_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(G113gat), .A3(new_n569_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  INV_X1    g682(.A(new_n879_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n885_), .ZN(G1340gat));
  INV_X1    g685(.A(G120gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n522_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n878_), .B(new_n888_), .C1(KEYINPUT60), .C2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n522_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n887_), .ZN(G1341gat));
  AOI21_X1  g690(.A(G127gat), .B1(new_n878_), .B2(new_n777_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n881_), .A2(G127gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n777_), .ZN(G1342gat));
  AOI21_X1  g693(.A(G134gat), .B1(new_n878_), .B2(new_n606_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n881_), .A2(G134gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n610_), .ZN(G1343gat));
  NOR3_X1   g696(.A1(new_n872_), .A2(new_n418_), .A3(new_n451_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(new_n668_), .A3(new_n424_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n752_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n213_), .ZN(G1344gat));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n522_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n214_), .ZN(G1345gat));
  NOR2_X1   g702(.A1(new_n899_), .A2(new_n635_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT61), .B(G155gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  NOR3_X1   g705(.A1(new_n899_), .A2(new_n588_), .A3(new_n675_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n899_), .A2(new_n839_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n588_), .B2(new_n908_), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n638_), .A2(new_n424_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n453_), .A2(new_n451_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n859_), .A2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n349_), .B1(new_n913_), .B2(new_n569_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT62), .Z(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n569_), .A3(new_n379_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1348gat));
  AOI21_X1  g716(.A(G176gat), .B1(new_n913_), .B2(new_n749_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n872_), .A2(new_n911_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n522_), .A2(new_n350_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1349gat));
  AOI21_X1  g720(.A(G183gat), .B1(new_n919_), .B2(new_n777_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n635_), .A2(new_n354_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n913_), .B2(new_n923_), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT125), .Z(G1350gat));
  INV_X1    g724(.A(new_n913_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G190gat), .B1(new_n926_), .B2(new_n675_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n606_), .A2(new_n355_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT126), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n926_), .B2(new_n929_), .ZN(G1351gat));
  NOR3_X1   g729(.A1(new_n872_), .A2(new_n453_), .A3(new_n451_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n910_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n752_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n525_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n522_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n237_), .A2(KEYINPUT127), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n237_), .A2(KEYINPUT127), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1353gat));
  NOR2_X1   g738(.A1(new_n932_), .A2(new_n635_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n940_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1354gat));
  INV_X1    g742(.A(new_n932_), .ZN(new_n944_));
  AOI21_X1  g743(.A(G218gat), .B1(new_n944_), .B2(new_n606_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n944_), .A2(G218gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n610_), .B2(new_n946_), .ZN(G1355gat));
endmodule


