//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OR3_X1    g006(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT65), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n211_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n208_), .A3(new_n210_), .A4(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT10), .B(G99gat), .Z(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT9), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(new_n225_), .A4(new_n207_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G43gat), .B(G50gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G36gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G29gat), .ZN(new_n230_));
  INV_X1    g029(.A(G29gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G36gat), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n230_), .A2(new_n232_), .A3(KEYINPUT71), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT71), .B1(new_n230_), .B2(new_n232_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n228_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n231_), .A2(G36gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n229_), .A2(G29gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n230_), .A2(new_n232_), .A3(KEYINPUT71), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n227_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n218_), .A2(KEYINPUT72), .A3(new_n226_), .A4(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT72), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n226_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n235_), .A2(new_n241_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(KEYINPUT68), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n250_), .B(new_n226_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n235_), .A2(new_n241_), .A3(KEYINPUT15), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT15), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT34), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n248_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G190gat), .B(G218gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT73), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G134gat), .B(G162gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT36), .ZN(new_n268_));
  INV_X1    g067(.A(new_n262_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n248_), .A2(new_n255_), .A3(new_n269_), .A4(new_n260_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n267_), .B(KEYINPUT36), .Z(new_n274_));
  AOI211_X1 g073(.A(new_n258_), .B(new_n259_), .C1(new_n248_), .C2(new_n255_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n270_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT75), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n279_), .B(new_n274_), .C1(new_n276_), .C2(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n202_), .B1(new_n273_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n271_), .B(KEYINPUT74), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT37), .A3(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G15gat), .B(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G1gat), .A2(G8gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT14), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n286_), .A2(new_n287_), .A3(new_n292_), .A4(new_n288_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G231gat), .A2(G233gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n300_));
  INV_X1    g099(.A(G64gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G57gat), .ZN(new_n302_));
  INV_X1    g101(.A(G57gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G64gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT11), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT67), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(new_n307_), .A3(KEYINPUT11), .ZN(new_n308_));
  XOR2_X1   g107(.A(G71gat), .B(G78gat), .Z(new_n309_));
  NAND4_X1  g108(.A1(new_n300_), .A2(new_n306_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(KEYINPUT11), .B2(new_n299_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n305_), .A2(KEYINPUT67), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n307_), .B1(new_n299_), .B2(KEYINPUT11), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n298_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n298_), .A2(new_n315_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G183gat), .B(G211gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT17), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT17), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n324_), .B1(new_n327_), .B2(new_n318_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n285_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT76), .ZN(new_n330_));
  INV_X1    g129(.A(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(G176gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT81), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(G169gat), .B2(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT25), .B(G183gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(G169gat), .B2(G176gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n338_), .A2(new_n343_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n350_), .A3(new_n342_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n341_), .A2(new_n350_), .A3(KEYINPUT82), .A4(new_n342_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n331_), .ZN(new_n356_));
  OAI21_X1  g155(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n349_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT30), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(G15gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT84), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G113gat), .B(G120gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT31), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n374_), .B2(KEYINPUT83), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n363_), .A2(new_n368_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n369_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n363_), .A2(new_n368_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n363_), .A2(new_n368_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n375_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n377_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G155gat), .ZN(new_n390_));
  INV_X1    g189(.A(G162gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT85), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(G155gat), .B2(G162gat), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n392_), .A2(new_n394_), .B1(G155gat), .B2(G162gat), .ZN(new_n395_));
  AND3_X1   g194(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  AND2_X1   g198(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT87), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n395_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G141gat), .B(G148gat), .Z(new_n410_));
  AND2_X1   g209(.A1(new_n392_), .A2(new_n394_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT1), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n410_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n373_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n373_), .A3(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT98), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n419_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n417_), .B2(KEYINPUT4), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(KEYINPUT4), .A3(new_n418_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT96), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n417_), .A2(new_n427_), .A3(KEYINPUT4), .A4(new_n418_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n424_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n389_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n424_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n409_), .A2(new_n373_), .A3(new_n414_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n373_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n427_), .B1(new_n434_), .B2(KEYINPUT4), .ZN(new_n435_));
  INV_X1    g234(.A(new_n428_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n420_), .B(KEYINPUT98), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n388_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n430_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n383_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT91), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT21), .ZN(new_n444_));
  INV_X1    g243(.A(G197gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G204gat), .ZN(new_n446_));
  INV_X1    g245(.A(G204gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G197gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G218gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G211gat), .ZN(new_n451_));
  INV_X1    g250(.A(G211gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G218gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n446_), .A2(new_n448_), .A3(KEYINPUT89), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n445_), .A3(G204gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT21), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G211gat), .B(G218gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n446_), .A2(new_n448_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(KEYINPUT21), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n455_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT90), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G197gat), .B(G204gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n454_), .B1(new_n444_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n446_), .A2(new_n448_), .A3(KEYINPUT89), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT21), .A3(new_n458_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n467_), .A2(new_n469_), .B1(new_n454_), .B2(new_n449_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G228gat), .A2(G233gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n465_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n443_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  AOI221_X4 g276(.A(KEYINPUT90), .B1(new_n454_), .B2(new_n449_), .C1(new_n467_), .C2(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n466_), .A2(new_n444_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n479_), .B(new_n461_), .C1(new_n456_), .C2(new_n459_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n471_), .B1(new_n480_), .B2(new_n455_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n476_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n482_), .A2(KEYINPUT91), .A3(new_n483_), .A4(new_n473_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n473_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n476_), .B2(new_n470_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT92), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n488_), .B(new_n485_), .C1(new_n476_), .C2(new_n470_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n477_), .A2(new_n484_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n442_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n409_), .A2(new_n475_), .A3(new_n414_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G22gat), .B(G50gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n495_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n477_), .A2(new_n484_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n487_), .A2(new_n489_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n504_), .A2(new_n492_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n492_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n493_), .A2(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n491_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n490_), .A2(new_n492_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n510_), .A2(new_n442_), .A3(new_n511_), .A4(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT27), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n349_), .A2(new_n359_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n356_), .A2(new_n357_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT95), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n351_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n343_), .A2(KEYINPUT95), .A3(new_n350_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n345_), .A2(KEYINPUT94), .ZN(new_n522_));
  INV_X1    g321(.A(G190gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT26), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT26), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(G190gat), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n524_), .A2(new_n526_), .A3(KEYINPUT94), .ZN(new_n527_));
  INV_X1    g326(.A(new_n344_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n522_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n338_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n521_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n464_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n516_), .A2(KEYINPUT20), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G226gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT19), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G8gat), .B(G36gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT18), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G64gat), .B(G92gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n338_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n345_), .A2(KEYINPUT94), .ZN(new_n544_));
  INV_X1    g343(.A(new_n527_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n344_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n543_), .A2(new_n546_), .B1(new_n520_), .B2(new_n519_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n542_), .B1(new_n547_), .B2(new_n470_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n535_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n465_), .A2(new_n472_), .A3(new_n360_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n536_), .A2(new_n541_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n541_), .B1(new_n536_), .B2(new_n551_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n514_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AND4_X1   g353(.A1(KEYINPUT20), .A2(new_n516_), .A3(new_n549_), .A4(new_n532_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n549_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n540_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n536_), .A2(new_n551_), .A3(new_n541_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(KEYINPUT27), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n513_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n441_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT100), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n508_), .A2(new_n512_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n430_), .A2(new_n439_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT33), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n439_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n552_), .A2(new_n553_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT33), .A4(new_n388_), .ZN(new_n571_));
  OAI221_X1 g370(.A(new_n419_), .B1(KEYINPUT4), .B2(new_n417_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n388_), .B1(new_n434_), .B2(new_n423_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n541_), .A2(KEYINPUT32), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT99), .B(new_n577_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n536_), .A2(new_n551_), .A3(new_n576_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n440_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n575_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n564_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n560_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n587_), .A2(new_n513_), .A3(KEYINPUT100), .A4(new_n565_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n567_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n562_), .B1(new_n589_), .B2(new_n383_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT12), .B1(new_n245_), .B2(new_n315_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n245_), .A2(new_n315_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n310_), .A2(new_n314_), .A3(KEYINPUT12), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n249_), .A2(new_n251_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n594_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n592_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n245_), .A2(new_n315_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n597_), .A2(new_n601_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n607_), .B(new_n609_), .C1(KEYINPUT69), .C2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n254_), .A2(new_n296_), .A3(new_n252_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n296_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(new_n242_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n242_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n296_), .B1(new_n241_), .B2(new_n235_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n625_), .A2(KEYINPUT77), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT78), .B(KEYINPUT79), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n625_), .B2(KEYINPUT77), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n621_), .A2(new_n624_), .A3(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT80), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT80), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n621_), .A2(new_n624_), .A3(new_n636_), .A4(new_n631_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n615_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n590_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n330_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n290_), .A3(new_n440_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n283_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n590_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n328_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n615_), .A4(new_n639_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G1gat), .B1(new_n650_), .B2(new_n565_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n644_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n651_), .A3(new_n652_), .ZN(G1324gat));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n291_), .A3(new_n560_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n650_), .A2(new_n587_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(KEYINPUT101), .A2(KEYINPUT39), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n291_), .B1(KEYINPUT101), .B2(KEYINPUT39), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT40), .B(new_n654_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(new_n383_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n642_), .A2(new_n365_), .A3(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT102), .ZN(new_n667_));
  OAI21_X1  g466(.A(G15gat), .B1(new_n650_), .B2(new_n383_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT41), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT41), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n667_), .A2(new_n669_), .A3(new_n670_), .ZN(G1326gat));
  OAI21_X1  g470(.A(G22gat), .B1(new_n650_), .B2(new_n564_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT42), .ZN(new_n673_));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n642_), .A2(new_n674_), .A3(new_n513_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1327gat));
  NOR2_X1   g475(.A1(new_n646_), .A2(new_n649_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT103), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n641_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n440_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n589_), .A2(new_n383_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n562_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n285_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n277_), .A2(KEYINPUT37), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n646_), .A2(new_n202_), .B1(new_n283_), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n590_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n640_), .A2(new_n649_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT44), .B1(new_n690_), .B2(new_n691_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n565_), .A2(new_n231_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n681_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n693_), .A2(new_n694_), .A3(new_n587_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n229_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n587_), .A2(KEYINPUT104), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n587_), .A2(KEYINPUT104), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n679_), .A2(G36gat), .A3(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n700_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n706_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n708_), .B(KEYINPUT46), .C1(new_n229_), .C2(new_n699_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1329gat));
  AOI21_X1  g509(.A(new_n685_), .B1(new_n684_), .B2(new_n285_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n590_), .A2(KEYINPUT43), .A3(new_n688_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n691_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n383_), .A2(new_n367_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n715_), .A2(KEYINPUT105), .A3(new_n692_), .A4(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n692_), .A3(new_n716_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G43gat), .B1(new_n680_), .B2(new_n665_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n723_));
  AND4_X1   g522(.A1(new_n717_), .A2(new_n720_), .A3(new_n722_), .A4(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n725_), .B2(new_n717_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n680_), .B2(new_n513_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n513_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n695_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1331gat));
  NOR3_X1   g531(.A1(new_n590_), .A2(new_n615_), .A3(new_n639_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n330_), .A2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(KEYINPUT108), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(KEYINPUT108), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n303_), .A3(new_n440_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n626_), .A2(new_n632_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n649_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n615_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n648_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n565_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n738_), .A2(new_n743_), .ZN(G1332gat));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n301_), .A3(new_n703_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G64gat), .B1(new_n742_), .B2(new_n704_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT48), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1333gat));
  NAND3_X1  g547(.A1(new_n648_), .A2(new_n665_), .A3(new_n741_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G71gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT109), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n752_), .A3(G71gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n383_), .A2(G71gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n735_), .A2(new_n736_), .A3(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n751_), .A2(KEYINPUT49), .A3(new_n753_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT110), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n756_), .A2(new_n758_), .A3(new_n762_), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n737_), .A2(new_n765_), .A3(new_n513_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G78gat), .B1(new_n742_), .B2(new_n564_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT50), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1335gat));
  NAND2_X1  g568(.A1(new_n733_), .A2(new_n678_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT111), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n223_), .A3(new_n440_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n615_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(new_n328_), .A3(new_n739_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n686_), .B2(new_n689_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n565_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(new_n777_), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n771_), .A2(new_n224_), .A3(new_n560_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G92gat), .B1(new_n776_), .B2(new_n704_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1337gat));
  AND2_X1   g580(.A1(new_n665_), .A2(new_n219_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n775_), .A2(new_n665_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n771_), .A2(new_n782_), .B1(G99gat), .B2(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n220_), .A3(new_n513_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n775_), .A2(new_n513_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(G106gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(G106gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n786_), .B(new_n792_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n622_), .A2(new_n623_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n618_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n623_), .A2(new_n617_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n631_), .B(new_n799_), .C1(new_n616_), .C2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n610_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n609_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT114), .B1(new_n739_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n639_), .A2(new_n807_), .A3(new_n609_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n593_), .A2(new_n596_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n598_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n597_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n593_), .A2(new_n596_), .A3(KEYINPUT55), .A4(new_n594_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n594_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n812_), .A2(new_n814_), .A3(new_n815_), .A4(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n606_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT116), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n809_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n819_), .B2(new_n606_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT56), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n804_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n797_), .B1(new_n827_), .B2(new_n647_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n826_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n806_), .B(new_n808_), .C1(new_n825_), .C2(KEYINPUT56), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n803_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT57), .A3(new_n646_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n820_), .A2(KEYINPUT56), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n819_), .A2(new_n822_), .A3(new_n606_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n802_), .A2(new_n609_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n834_), .A4(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT117), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n835_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n834_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n802_), .A2(new_n609_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n820_), .B2(KEYINPUT56), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(KEYINPUT58), .A4(new_n834_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n837_), .A2(new_n841_), .A3(new_n285_), .A4(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n828_), .A2(new_n832_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n328_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n740_), .A2(KEYINPUT113), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n639_), .A2(new_n328_), .A3(KEYINPUT113), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n850_), .A2(new_n615_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n688_), .B2(new_n852_), .ZN(new_n853_));
  AND4_X1   g652(.A1(new_n849_), .A2(new_n852_), .A3(new_n282_), .A4(new_n284_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n848_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n561_), .A2(new_n665_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n440_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n639_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n855_), .B1(new_n847_), .B2(new_n328_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n565_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT59), .A3(new_n859_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n739_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n863_), .B1(new_n869_), .B2(new_n862_), .ZN(G1340gat));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n615_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n861_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n615_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n871_), .ZN(G1341gat));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877_));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n328_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n860_), .B2(new_n328_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n876_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n880_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT59), .B1(new_n867_), .B2(new_n859_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n866_), .A2(new_n864_), .A3(new_n565_), .A4(new_n858_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(KEYINPUT119), .A3(new_n882_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n884_), .A2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n861_), .B2(new_n647_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n865_), .A2(new_n868_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT120), .B(G134gat), .Z(new_n893_));
  NOR2_X1   g692(.A1(new_n688_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n892_), .B2(new_n894_), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n857_), .A2(new_n440_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n703_), .A2(new_n665_), .A3(new_n564_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n639_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n773_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n649_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  NAND4_X1  g705(.A1(new_n867_), .A2(new_n391_), .A3(new_n647_), .A4(new_n897_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n896_), .A2(new_n688_), .A3(new_n898_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n391_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT121), .B(new_n907_), .C1(new_n908_), .C2(new_n391_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1347gat));
  NAND3_X1  g712(.A1(new_n703_), .A2(new_n564_), .A3(new_n441_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT22), .B(G169gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n639_), .A3(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n918_));
  INV_X1    g717(.A(new_n914_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n857_), .A2(new_n639_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n915_), .A2(KEYINPUT122), .A3(new_n639_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n331_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n918_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(KEYINPUT122), .B1(new_n915_), .B2(new_n639_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n866_), .A2(new_n921_), .A3(new_n739_), .A4(new_n914_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n918_), .B(new_n925_), .C1(new_n927_), .C2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n917_), .B1(new_n926_), .B2(new_n930_), .ZN(G1348gat));
  NAND2_X1  g730(.A1(new_n915_), .A2(new_n773_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g732(.A1(new_n915_), .A2(new_n649_), .ZN(new_n934_));
  MUX2_X1   g733(.A(new_n344_), .B(G183gat), .S(new_n934_), .Z(G1350gat));
  INV_X1    g734(.A(new_n915_), .ZN(new_n936_));
  OAI21_X1  g735(.A(G190gat), .B1(new_n936_), .B2(new_n688_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n647_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n936_), .B2(new_n938_), .ZN(G1351gat));
  NAND3_X1  g738(.A1(new_n383_), .A2(new_n513_), .A3(new_n565_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n866_), .A2(new_n704_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n639_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n942_), .B2(new_n445_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n445_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n941_), .A2(new_n945_), .A3(G197gat), .A4(new_n639_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n943_), .A2(new_n944_), .A3(new_n946_), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n941_), .A2(new_n773_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n447_), .A2(KEYINPUT125), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT126), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n948_), .B(new_n950_), .ZN(G1353gat));
  AOI21_X1  g750(.A(new_n328_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT127), .Z(new_n953_));
  NAND2_X1  g752(.A1(new_n941_), .A2(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n954_), .B(new_n955_), .Z(G1354gat));
  NAND3_X1  g755(.A1(new_n941_), .A2(new_n450_), .A3(new_n647_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n941_), .A2(new_n285_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n450_), .ZN(G1355gat));
endmodule


