//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n203_), .A2(new_n204_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n211_));
  OAI22_X1  g010(.A1(new_n210_), .A2(new_n211_), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT6), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT65), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(new_n218_), .B2(new_n220_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n212_), .B(new_n216_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n225_));
  OR2_X1    g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT68), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n225_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n218_), .A2(new_n220_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n212_), .A2(new_n234_), .A3(new_n216_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n224_), .A2(new_n233_), .B1(new_n237_), .B2(KEYINPUT8), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n222_), .A2(new_n223_), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n240_), .B(new_n230_), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n226_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n228_), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n215_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n239_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n209_), .B1(new_n238_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n239_), .A2(new_n246_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n208_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n225_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n236_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n223_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n221_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n212_), .A2(new_n216_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT8), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n249_), .B(new_n251_), .C1(new_n257_), .C2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n248_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n260_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n249_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT12), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n209_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G176gat), .B(G204gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n270_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT69), .B(new_n275_), .C1(new_n263_), .C2(new_n269_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT13), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT13), .B1(new_n277_), .B2(new_n278_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT70), .ZN(new_n283_));
  INV_X1    g082(.A(new_n281_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n279_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(KEYINPUT71), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(KEYINPUT71), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT34), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n238_), .A2(new_n247_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G29gat), .B(G36gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n296_), .B(KEYINPUT72), .ZN(new_n301_));
  INV_X1    g100(.A(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n301_), .A2(new_n302_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n298_), .A2(new_n299_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n295_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n266_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT35), .B(new_n294_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n305_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n266_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n294_), .A2(KEYINPUT35), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n307_), .A2(new_n308_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n295_), .A2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n294_), .A2(KEYINPUT35), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G190gat), .B(G218gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(G134gat), .B(G162gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n312_), .A2(new_n319_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT77), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n312_), .A2(new_n329_), .A3(new_n319_), .A4(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n324_), .B(KEYINPUT36), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT37), .B1(new_n331_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT37), .ZN(new_n337_));
  AOI211_X1 g136(.A(new_n337_), .B(new_n334_), .C1(new_n328_), .C2(new_n330_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G155gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G183gat), .B(G211gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G1gat), .ZN(new_n348_));
  INV_X1    g147(.A(G8gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT14), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G15gat), .ZN(new_n351_));
  INV_X1    g150(.A(G22gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G15gat), .A2(G22gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT79), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n356_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G1gat), .B(G8gat), .Z(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n366_));
  OAI211_X1 g165(.A(G231gat), .B(G233gat), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G231gat), .A2(G233gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n251_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n251_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n373_));
  OAI221_X1 g172(.A(new_n347_), .B1(KEYINPUT17), .B2(new_n345_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n372_), .A2(new_n347_), .A3(new_n373_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n340_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n292_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT82), .Z(new_n379_));
  INV_X1    g178(.A(G169gat), .ZN(new_n380_));
  INV_X1    g179(.A(G176gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT24), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT25), .B(G183gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT26), .B(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n382_), .A2(KEYINPUT84), .A3(KEYINPUT24), .A4(new_n383_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT85), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n386_), .A2(new_n389_), .A3(new_n393_), .A4(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n395_), .B(KEYINPUT86), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n397_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n382_), .A2(KEYINPUT24), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n392_), .A2(new_n394_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n396_), .A2(KEYINPUT23), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n399_), .B2(KEYINPUT23), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n403_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(G71gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(G99gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n413_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G127gat), .B(G134gat), .Z(new_n419_));
  XOR2_X1   g218(.A(G113gat), .B(G120gat), .Z(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n418_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G15gat), .B(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT87), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT30), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT31), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n422_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G85gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT0), .B(G57gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(KEYINPUT1), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(KEYINPUT1), .B2(new_n433_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n421_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n439_), .B(KEYINPUT2), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT3), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n437_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n437_), .A2(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT3), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n442_), .A2(new_n447_), .A3(KEYINPUT89), .A4(new_n445_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n434_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n433_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n440_), .B(new_n441_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n440_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n421_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(KEYINPUT4), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n455_), .A2(new_n458_), .A3(KEYINPUT92), .A4(KEYINPUT4), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(new_n458_), .B2(KEYINPUT4), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n455_), .A2(new_n458_), .A3(new_n465_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(new_n464_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n432_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n472_), .A2(new_n464_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n470_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n472_), .B2(new_n464_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n477_), .A3(new_n431_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n427_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n456_), .A2(new_n457_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT29), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT28), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G22gat), .B(G50gat), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  INV_X1    g285(.A(G204gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(G197gat), .ZN(new_n488_));
  INV_X1    g287(.A(G197gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(G204gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT21), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G211gat), .B(G218gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(KEYINPUT91), .B2(new_n488_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n491_), .B(new_n492_), .C1(new_n495_), .C2(KEYINPUT21), .ZN(new_n496_));
  INV_X1    g295(.A(new_n492_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(KEYINPUT21), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT90), .B(new_n499_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G228gat), .A2(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(G78gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n215_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(new_n504_), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n485_), .A2(new_n486_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n413_), .A2(new_n499_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n405_), .B1(new_n400_), .B2(new_n409_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n408_), .A2(new_n384_), .A3(new_n389_), .A4(new_n402_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n496_), .A2(new_n498_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(KEYINPUT20), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT19), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n403_), .A3(new_n412_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n511_), .A2(new_n512_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n523_), .B2(new_n499_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n524_), .A3(new_n518_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G8gat), .B(G36gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT18), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G64gat), .B(G92gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n520_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n522_), .B1(new_n413_), .B2(new_n499_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n518_), .B1(new_n532_), .B2(new_n515_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n525_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n529_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n531_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(KEYINPUT96), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n529_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n499_), .B1(new_n523_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n541_), .B2(new_n523_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n519_), .B1(new_n543_), .B2(new_n532_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n521_), .A2(new_n524_), .A3(new_n519_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n530_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n538_), .A2(new_n540_), .A3(new_n546_), .ZN(new_n547_));
  AOI211_X1 g346(.A(KEYINPUT97), .B(new_n537_), .C1(KEYINPUT27), .C2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(KEYINPUT27), .ZN(new_n550_));
  INV_X1    g349(.A(new_n537_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n479_), .B(new_n509_), .C1(new_n548_), .C2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n478_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n475_), .A2(new_n477_), .A3(new_n431_), .A4(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n455_), .A2(new_n458_), .A3(new_n466_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n461_), .A2(new_n462_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n465_), .B1(new_n458_), .B2(KEYINPUT4), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n432_), .B(new_n558_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n561_), .A2(new_n535_), .A3(new_n531_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n544_), .A2(new_n545_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n533_), .A2(new_n534_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n529_), .A2(KEYINPUT32), .ZN(new_n566_));
  MUX2_X1   g365(.A(new_n564_), .B(new_n565_), .S(new_n566_), .Z(new_n567_));
  NOR3_X1   g366(.A1(new_n471_), .A2(new_n432_), .A3(new_n473_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n431_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n563_), .A2(new_n509_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n474_), .A2(new_n478_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n537_), .B1(new_n547_), .B2(KEYINPUT27), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n508_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n427_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n553_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n313_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n368_), .A2(new_n364_), .A3(new_n316_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  OAI22_X1  g380(.A1(new_n365_), .A2(new_n366_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n582_), .B2(new_n579_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT83), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G169gat), .B(G197gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(KEYINPUT83), .B(new_n587_), .C1(new_n581_), .C2(new_n583_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n577_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT98), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n379_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n348_), .A3(new_n572_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n594_), .A2(KEYINPUT38), .A3(new_n348_), .A4(new_n572_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n331_), .A2(new_n335_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT99), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n563_), .A2(new_n509_), .A3(new_n570_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n575_), .A3(new_n574_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n602_), .B2(new_n553_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n376_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n591_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n288_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n572_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n597_), .A2(new_n598_), .A3(new_n610_), .ZN(G1324gat));
  OR2_X1    g410(.A1(new_n548_), .A2(new_n552_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n379_), .A2(new_n349_), .A3(new_n613_), .A4(new_n593_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n607_), .A2(new_n613_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n616_), .B2(G8gat), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n615_), .A3(G8gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1325gat));
  NAND3_X1  g424(.A1(new_n594_), .A2(new_n351_), .A3(new_n427_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n351_), .B1(new_n607_), .B2(new_n427_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT41), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1326gat));
  XNOR2_X1  g428(.A(new_n508_), .B(KEYINPUT101), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n594_), .A2(new_n352_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n352_), .B1(new_n607_), .B2(new_n631_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT42), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1327gat));
  NAND2_X1  g434(.A1(new_n600_), .A2(new_n376_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n288_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n593_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n638_), .B2(new_n572_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n283_), .A2(new_n287_), .A3(new_n591_), .A4(new_n376_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n339_), .B(KEYINPUT103), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n577_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n340_), .A2(new_n643_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n602_), .B2(new_n553_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT44), .B(new_n642_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n572_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n639_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  NOR2_X1   g453(.A1(new_n612_), .A2(G36gat), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n592_), .A2(KEYINPUT98), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n592_), .A2(KEYINPUT98), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n637_), .B(new_n655_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT45), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n650_), .A2(new_n613_), .A3(new_n651_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT104), .B1(new_n660_), .B2(G36gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n660_), .A2(G36gat), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n660_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n673_), .A2(new_n664_), .A3(new_n665_), .A4(new_n659_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n668_), .A2(new_n674_), .ZN(G1329gat));
  AOI21_X1  g474(.A(G43gat), .B1(new_n638_), .B2(new_n427_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n427_), .A2(G43gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n652_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1330gat));
  INV_X1    g479(.A(G50gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n638_), .A2(new_n681_), .A3(new_n631_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n652_), .A2(new_n508_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(new_n681_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT106), .ZN(G1331gat));
  NAND2_X1  g484(.A1(new_n577_), .A2(new_n605_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT107), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(new_n377_), .A3(new_n288_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n688_), .A2(KEYINPUT108), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(KEYINPUT108), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n572_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(G57gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n591_), .A2(new_n376_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n291_), .A2(new_n603_), .A3(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n609_), .A2(new_n692_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n691_), .A2(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(G1332gat));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n694_), .B2(new_n613_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT48), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(new_n697_), .A3(new_n613_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1333gat));
  NAND2_X1  g500(.A1(new_n694_), .A2(new_n427_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(G71gat), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT49), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n702_), .B2(G71gat), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n688_), .A2(new_n415_), .A3(new_n427_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(G1334gat));
  AOI21_X1  g510(.A(new_n502_), .B1(new_n694_), .B2(new_n631_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT50), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n688_), .A2(new_n502_), .A3(new_n631_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n292_), .A2(new_n636_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n687_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G85gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n572_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n645_), .A2(new_n647_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n288_), .A2(new_n605_), .A3(new_n376_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n721_), .A2(new_n609_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n719_), .B2(new_n723_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n718_), .B2(new_n613_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n721_), .A2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n613_), .A2(G92gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT110), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n726_), .B2(new_n728_), .ZN(G1337gat));
  AOI21_X1  g528(.A(new_n214_), .B1(new_n726_), .B2(new_n427_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n427_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n718_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n726_), .A2(new_n508_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G106gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT52), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n718_), .A2(new_n215_), .A3(new_n508_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(KEYINPUT52), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n735_), .B2(G106gat), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n738_), .B(new_n734_), .C1(new_n740_), .C2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n739_), .A2(new_n744_), .ZN(G1339gat));
  NAND3_X1  g544(.A1(new_n339_), .A2(new_n282_), .A3(new_n693_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT54), .B1(new_n746_), .B2(KEYINPUT112), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n282_), .A2(new_n693_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .A4(new_n339_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n339_), .A2(new_n749_), .A3(new_n282_), .A4(new_n693_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n747_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n747_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n757_));
  INV_X1    g556(.A(new_n580_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n578_), .A2(new_n579_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n582_), .B2(new_n579_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n588_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n587_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n278_), .A2(new_n277_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n269_), .A2(KEYINPUT55), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n265_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n265_), .A2(new_n268_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT55), .B1(new_n766_), .B2(new_n262_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n764_), .B(new_n765_), .C1(new_n767_), .C2(KEYINPUT114), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n269_), .A2(new_n769_), .A3(KEYINPUT55), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n275_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n766_), .A2(new_n262_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT114), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n769_), .B1(new_n269_), .B2(KEYINPUT55), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n764_), .A4(new_n765_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n773_), .A2(new_n774_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n270_), .A2(new_n276_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n589_), .A2(new_n590_), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n275_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(KEYINPUT115), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n763_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n757_), .B1(new_n786_), .B2(new_n600_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n787_), .A2(KEYINPUT117), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n600_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(KEYINPUT117), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n761_), .A2(new_n762_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n780_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n784_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n793_), .B(KEYINPUT58), .C1(new_n794_), .C2(new_n784_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n340_), .A3(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n788_), .A2(new_n791_), .A3(new_n792_), .A4(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n756_), .B1(new_n800_), .B2(new_n376_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n612_), .A2(new_n509_), .A3(new_n572_), .A4(new_n427_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n802_), .A2(KEYINPUT118), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(KEYINPUT118), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n801_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT119), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(KEYINPUT59), .C1(new_n801_), .C2(new_n805_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n787_), .A2(new_n799_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n790_), .B1(new_n813_), .B2(KEYINPUT120), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n787_), .A2(new_n815_), .A3(new_n799_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n604_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n756_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n805_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n807_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n812_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n754_), .A2(new_n755_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n787_), .A2(new_n815_), .A3(new_n799_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n815_), .B1(new_n787_), .B2(new_n799_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n790_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n822_), .B1(new_n825_), .B2(new_n604_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n807_), .A4(new_n819_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n811_), .A2(new_n591_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G113gat), .ZN(new_n830_));
  INV_X1    g629(.A(new_n806_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n831_), .A2(G113gat), .A3(new_n605_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1340gat));
  NAND3_X1  g632(.A1(new_n811_), .A2(new_n291_), .A3(new_n828_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT122), .B(G120gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n288_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n838_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(KEYINPUT60), .B2(new_n835_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n831_), .A2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT123), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n837_), .A2(new_n842_), .ZN(G1341gat));
  NAND3_X1  g642(.A1(new_n811_), .A2(new_n604_), .A3(new_n828_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G127gat), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n831_), .A2(G127gat), .A3(new_n376_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1342gat));
  NAND3_X1  g646(.A1(new_n811_), .A2(new_n340_), .A3(new_n828_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G134gat), .ZN(new_n849_));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n806_), .A2(new_n850_), .A3(new_n600_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n800_), .A2(new_n376_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n822_), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n613_), .A2(new_n509_), .A3(new_n609_), .A4(new_n427_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n591_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT124), .B(G141gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n291_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n604_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  AOI21_X1  g663(.A(G162gat), .B1(new_n856_), .B2(new_n600_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n644_), .A2(G162gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n856_), .B2(new_n866_), .ZN(G1347gat));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n612_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n630_), .B(new_n869_), .C1(new_n817_), .C2(new_n756_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n605_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT22), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G169gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n380_), .B1(new_n871_), .B2(new_n868_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n875_), .ZN(G1348gat));
  NAND2_X1  g675(.A1(new_n854_), .A2(new_n509_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n291_), .A2(G176gat), .A3(new_n869_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n870_), .A2(new_n838_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n381_), .B2(new_n880_), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n869_), .A2(new_n604_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n877_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G183gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n818_), .A2(new_n631_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n387_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1350gat));
  NAND4_X1  g686(.A1(new_n885_), .A2(new_n388_), .A3(new_n600_), .A4(new_n869_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(G190gat), .C1(new_n870_), .C2(new_n339_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n826_), .A2(new_n340_), .A3(new_n630_), .A4(new_n869_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n892_), .B2(G190gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n888_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n896_), .B(new_n888_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1351gat));
  NAND3_X1  g697(.A1(new_n609_), .A2(new_n508_), .A3(new_n575_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n801_), .A2(new_n612_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n591_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n291_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n604_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT63), .B(G211gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908_));
  INV_X1    g707(.A(G211gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n905_), .A2(KEYINPUT127), .A3(new_n908_), .A4(new_n909_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n907_), .B1(new_n912_), .B2(new_n913_), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n900_), .A2(new_n915_), .A3(new_n600_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n900_), .A2(new_n340_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n915_), .ZN(G1355gat));
endmodule


