//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT13), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G71gat), .B(G78gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(KEYINPUT11), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT68), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(KEYINPUT11), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT66), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n217_), .A2(new_n222_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n216_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT7), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT6), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n221_), .A2(new_n223_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  AND2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n220_), .A2(KEYINPUT66), .B1(KEYINPUT7), .B2(new_n224_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n226_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT67), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n234_), .A2(new_n223_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n240_), .A2(new_n232_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n233_), .B1(new_n241_), .B2(new_n229_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(G92gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G85gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(KEYINPUT9), .B2(new_n230_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT10), .B(G99gat), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n216_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n227_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n213_), .A2(new_n242_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n211_), .B(new_n212_), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT12), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n229_), .B1(new_n240_), .B2(new_n232_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n250_), .B(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n253_), .B1(new_n257_), .B2(new_n250_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G230gat), .ZN(new_n265_));
  INV_X1    g064(.A(G233gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n252_), .A2(KEYINPUT69), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n252_), .A2(KEYINPUT69), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n263_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G120gat), .B(G148gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n279_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n269_), .A2(new_n273_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n207_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n282_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n284_), .B(new_n285_), .C1(new_n286_), .C2(new_n205_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n205_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n288_), .B2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT78), .B(G1gat), .Z(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G43gat), .B(G50gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G229gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT80), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT81), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT81), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n297_), .B(new_n301_), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G229gat), .A3(G233gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G141gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G169gat), .B(G197gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n316_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n290_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT99), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT99), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n290_), .A2(new_n322_), .A3(new_n319_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  XNOR2_X1  g126(.A(G141gat), .B(G148gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT1), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n331_), .B2(KEYINPUT1), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(G155gat), .B2(G162gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT85), .A3(new_n329_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n328_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n329_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(new_n331_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342_));
  INV_X1    g141(.A(G141gat), .ZN(new_n343_));
  INV_X1    g142(.A(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n345_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT86), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n341_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n327_), .B1(new_n338_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT86), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n352_), .B(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n340_), .B1(new_n357_), .B2(new_n350_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n325_), .B(new_n326_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n336_), .A2(KEYINPUT85), .A3(new_n329_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT85), .B1(new_n336_), .B2(new_n329_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n330_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n358_), .B(new_n359_), .C1(new_n362_), .C2(new_n328_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n355_), .A2(new_n363_), .A3(KEYINPUT4), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT93), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n355_), .A2(new_n363_), .A3(new_n366_), .A4(KEYINPUT4), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT94), .Z(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n355_), .B2(KEYINPUT4), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n355_), .A2(new_n363_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G85gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT0), .B(G57gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  NAND3_X1  g179(.A1(new_n373_), .A2(new_n376_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n382_));
  INV_X1    g181(.A(new_n380_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n371_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n376_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n381_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  NOR3_X1   g191(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT24), .ZN(new_n395_));
  INV_X1    g194(.A(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G183gat), .ZN(new_n402_));
  INV_X1    g201(.A(G183gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT25), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G190gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT23), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(G183gat), .A3(G190gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT84), .B(KEYINPUT23), .C1(new_n403_), .C2(new_n406_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n399_), .A2(new_n405_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n403_), .A2(new_n406_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n394_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT22), .B(G169gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n397_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI211_X1 g220(.A(KEYINPUT92), .B(new_n417_), .C1(new_n418_), .C2(new_n397_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n413_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT21), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G197gat), .A2(G204gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G197gat), .A2(G204gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(G204gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(KEYINPUT21), .A3(new_n425_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G211gat), .B(G218gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT88), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n428_), .A2(new_n432_), .A3(new_n436_), .A4(new_n433_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n432_), .A2(new_n433_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n423_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n438_), .B1(new_n434_), .B2(KEYINPUT88), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT89), .A3(new_n437_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n402_), .A2(new_n404_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT82), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n403_), .B2(KEYINPUT25), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(KEYINPUT83), .A3(new_n400_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n400_), .A2(new_n450_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n399_), .A2(new_n414_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n411_), .A2(new_n415_), .A3(new_n412_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n456_), .A2(new_n457_), .B1(new_n419_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n441_), .B1(new_n446_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT20), .B1(new_n423_), .B2(new_n440_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT95), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n392_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  AND4_X1   g263(.A1(KEYINPUT89), .A2(new_n435_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT89), .B1(new_n444_), .B2(new_n437_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n459_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n392_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n423_), .B2(new_n440_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n464_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G8gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT18), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G64gat), .B(G92gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n467_), .A2(new_n470_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n392_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n476_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n407_), .A2(new_n410_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT22), .B(G169gat), .Z(new_n482_));
  OAI21_X1  g281(.A(new_n394_), .B1(new_n482_), .B2(G176gat), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n483_), .B2(KEYINPUT92), .ZN(new_n484_));
  INV_X1    g283(.A(new_n422_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n399_), .A2(new_n405_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n411_), .A2(new_n412_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n484_), .A2(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n440_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n469_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n490_), .B(new_n468_), .C1(new_n446_), .C2(new_n459_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n479_), .A2(new_n480_), .A3(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n477_), .A2(KEYINPUT98), .A3(KEYINPUT27), .A4(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n468_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT20), .B(new_n468_), .C1(new_n423_), .C2(new_n440_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n465_), .A2(new_n466_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n459_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n476_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT27), .B1(new_n492_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT98), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n492_), .A2(KEYINPUT27), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n480_), .B1(new_n464_), .B2(new_n471_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n493_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G22gat), .B(G50gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n338_), .A2(new_n354_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n508_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n512_), .A3(new_n507_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n515_), .A2(new_n517_), .A3(KEYINPUT91), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT91), .B1(new_n515_), .B2(new_n517_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(G228gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(G228gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n266_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT29), .B1(new_n338_), .B2(new_n354_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n496_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G78gat), .B(G106gat), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n489_), .B1(KEYINPUT90), .B2(new_n527_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n532_), .B(KEYINPUT29), .C1(new_n338_), .C2(new_n354_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n528_), .B(new_n530_), .C1(new_n534_), .C2(new_n526_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n528_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n526_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n520_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(new_n518_), .A3(new_n538_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G71gat), .B(G99gat), .ZN(new_n543_));
  INV_X1    g342(.A(G43gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n459_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n359_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G227gat), .A2(G233gat), .ZN(new_n548_));
  INV_X1    g347(.A(G15gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT30), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT31), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n547_), .A2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR4_X1   g355(.A1(new_n390_), .A2(new_n506_), .A3(new_n542_), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n383_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n373_), .A2(new_n376_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n380_), .B1(new_n374_), .B2(new_n370_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n365_), .A2(new_n367_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n375_), .B1(new_n355_), .B2(KEYINPUT4), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  AND4_X1   g363(.A1(new_n492_), .A2(new_n560_), .A3(new_n564_), .A4(new_n499_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n381_), .A2(new_n558_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n381_), .A2(new_n386_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n494_), .A2(new_n498_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n472_), .B2(new_n568_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n565_), .A2(new_n566_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT96), .B1(new_n571_), .B2(new_n542_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n477_), .A2(KEYINPUT27), .A3(new_n492_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n500_), .B1(new_n573_), .B2(new_n502_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n574_), .A2(new_n389_), .A3(new_n542_), .A4(new_n493_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n492_), .A2(new_n499_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(new_n566_), .A3(new_n560_), .A4(new_n564_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n472_), .A2(new_n568_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n569_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n567_), .A3(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n577_), .A2(new_n580_), .B1(new_n541_), .B2(new_n540_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n572_), .A2(new_n575_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n557_), .B1(new_n584_), .B2(new_n556_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT36), .Z(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT34), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n301_), .B(new_n251_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n303_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n595_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n303_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n250_), .B(KEYINPUT70), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n242_), .B2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n604_), .A2(new_n598_), .A3(new_n594_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n589_), .B1(new_n601_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n594_), .B1(new_n604_), .B2(new_n598_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT100), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n585_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n213_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n298_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n617_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n617_), .A2(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n324_), .A2(new_n614_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n202_), .B1(new_n630_), .B2(new_n390_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT101), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT74), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n290_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n287_), .A2(new_n289_), .A3(KEYINPUT74), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT37), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n606_), .A2(new_n637_), .A3(new_n610_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT77), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(KEYINPUT77), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT76), .ZN(new_n642_));
  INV_X1    g441(.A(new_n589_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT75), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n610_), .B1(new_n644_), .B2(KEYINPUT75), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n642_), .B(KEYINPUT37), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT75), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n606_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n610_), .A3(new_n645_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n642_), .B1(new_n652_), .B2(KEYINPUT37), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n641_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n628_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n636_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n319_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n585_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(new_n390_), .A3(new_n291_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n632_), .A2(new_n663_), .A3(new_n664_), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n630_), .A2(new_n506_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G8gat), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n506_), .A2(new_n292_), .ZN(new_n670_));
  OAI22_X1  g469(.A1(new_n668_), .A2(new_n669_), .B1(new_n660_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI221_X1 g472(.A(KEYINPUT40), .B1(new_n660_), .B2(new_n670_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  INV_X1    g474(.A(new_n556_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n549_), .B1(new_n630_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n661_), .A2(new_n549_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n678_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  INV_X1    g481(.A(G22gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n630_), .B2(new_n542_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT42), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n661_), .A2(new_n683_), .A3(new_n542_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1327gat));
  NAND3_X1  g486(.A1(new_n321_), .A2(new_n628_), .A3(new_n323_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n540_), .B(new_n541_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n691_));
  OAI22_X1  g490(.A1(new_n581_), .A2(new_n582_), .B1(new_n506_), .B2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n571_), .A2(new_n542_), .A3(KEYINPUT96), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n556_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n557_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n655_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT104), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n585_), .B2(new_n654_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n696_), .A2(new_n701_), .A3(new_n697_), .A4(new_n655_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n390_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n690_), .B2(new_n703_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G29gat), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n629_), .A2(new_n612_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n290_), .A2(new_n659_), .A3(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT105), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n389_), .A2(G29gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT106), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n707_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n707_), .A2(KEYINPUT107), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1328gat));
  NAND2_X1  g517(.A1(new_n704_), .A2(new_n506_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G36gat), .B1(new_n719_), .B2(new_n706_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n721_));
  NOR2_X1   g520(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n722_));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n710_), .A2(new_n723_), .A3(new_n506_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n725_));
  OR2_X1    g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n725_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n722_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n720_), .A2(new_n721_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n721_), .B1(new_n720_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  INV_X1    g530(.A(new_n710_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n544_), .B1(new_n732_), .B2(new_n556_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n704_), .A2(G43gat), .A3(new_n676_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n706_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g535(.A1(new_n704_), .A2(new_n542_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G50gat), .B1(new_n737_), .B2(new_n706_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n542_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(G50gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT111), .Z(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n732_), .B2(new_n741_), .ZN(G1331gat));
  NOR2_X1   g541(.A1(new_n319_), .A2(new_n628_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n634_), .A2(new_n614_), .A3(new_n635_), .A4(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n389_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n290_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n585_), .A2(new_n319_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n656_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G57gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n390_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n745_), .A2(new_n750_), .ZN(G1332gat));
  INV_X1    g550(.A(G64gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n752_), .A3(new_n506_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n506_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n744_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(G64gat), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(G1333gat));
  INV_X1    g558(.A(G71gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n748_), .A2(new_n760_), .A3(new_n676_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G71gat), .B1(new_n744_), .B2(new_n556_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT49), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT49), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1334gat));
  NOR2_X1   g564(.A1(new_n739_), .A2(G78gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT113), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n748_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G78gat), .B1(new_n744_), .B2(new_n739_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  NAND3_X1  g571(.A1(new_n746_), .A2(new_n628_), .A3(new_n658_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n702_), .A2(new_n700_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n654_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n701_), .B1(new_n775_), .B2(new_n697_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT114), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n699_), .A2(new_n778_), .A3(new_n700_), .A4(new_n702_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n773_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n389_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n634_), .A2(new_n635_), .A3(new_n708_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n747_), .ZN(new_n784_));
  INV_X1    g583(.A(G85gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n390_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(G1336gat));
  AOI21_X1  g586(.A(G92gat), .B1(new_n784_), .B2(new_n506_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n506_), .A2(new_n243_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n780_), .B2(new_n789_), .ZN(G1337gat));
  AOI21_X1  g589(.A(new_n215_), .B1(new_n780_), .B2(new_n676_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n783_), .A2(new_n676_), .A3(new_n247_), .A4(new_n747_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT115), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n556_), .B(new_n773_), .C1(new_n777_), .C2(new_n779_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n795_), .B(new_n792_), .C1(new_n796_), .C2(new_n215_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(KEYINPUT51), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n780_), .A2(new_n676_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n793_), .B1(new_n800_), .B2(G99gat), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n794_), .A2(new_n799_), .A3(KEYINPUT51), .A4(new_n797_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1338gat));
  NOR2_X1   g608(.A1(new_n773_), .A2(new_n739_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n216_), .B1(new_n810_), .B2(new_n703_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n784_), .A2(new_n216_), .A3(new_n542_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g615(.A(new_n743_), .B1(new_n288_), .B2(new_n283_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n655_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n817_), .B2(new_n655_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(KEYINPUT54), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n818_), .B(new_n822_), .C1(new_n817_), .C2(new_n655_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n311_), .A2(new_n307_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n305_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n825_), .B(new_n316_), .C1(new_n826_), .C2(new_n307_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n317_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n282_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT55), .B1(new_n264_), .B2(new_n268_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n269_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n264_), .A2(KEYINPUT55), .A3(new_n268_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n281_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT56), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n829_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n834_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(KEYINPUT56), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT120), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n836_), .A2(KEYINPUT58), .A3(new_n839_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n655_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n838_), .A2(KEYINPUT119), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n319_), .A2(new_n282_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n837_), .A2(KEYINPUT119), .A3(new_n838_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n848_), .A2(new_n849_), .B1(new_n286_), .B2(new_n828_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n613_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n849_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n828_), .A2(new_n286_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n844_), .A2(new_n851_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n824_), .B1(new_n856_), .B2(new_n628_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n506_), .A2(new_n542_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n390_), .A3(new_n676_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n319_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n628_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n824_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n859_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(KEYINPUT59), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n658_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n862_), .B1(new_n870_), .B2(new_n861_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n862_), .B(KEYINPUT121), .C1(new_n870_), .C2(new_n861_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1340gat));
  NOR2_X1   g674(.A1(new_n290_), .A2(KEYINPUT60), .ZN(new_n876_));
  MUX2_X1   g675(.A(new_n876_), .B(KEYINPUT60), .S(G120gat), .Z(new_n877_));
  NAND2_X1  g676(.A1(new_n860_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n636_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G120gat), .B1(new_n879_), .B2(new_n880_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n881_), .B2(new_n882_), .ZN(G1341gat));
  AOI21_X1  g682(.A(G127gat), .B1(new_n860_), .B2(new_n629_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n884_), .A2(KEYINPUT123), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(KEYINPUT123), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n867_), .A2(new_n869_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n629_), .A2(G127gat), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n860_), .A2(new_n890_), .A3(new_n613_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n654_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n890_), .ZN(G1343gat));
  NOR3_X1   g692(.A1(new_n857_), .A2(new_n739_), .A3(new_n676_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n506_), .A2(new_n389_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n658_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n343_), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n636_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n344_), .ZN(G1345gat));
  NOR2_X1   g699(.A1(new_n896_), .A2(new_n628_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT61), .B(G155gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n896_), .A2(new_n904_), .A3(new_n654_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n896_), .B2(new_n612_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT124), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n908_), .B(new_n904_), .C1(new_n896_), .C2(new_n612_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n905_), .B1(new_n907_), .B2(new_n909_), .ZN(G1347gat));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n396_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n390_), .A2(new_n556_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(new_n739_), .A3(new_n506_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n857_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n913_), .B1(new_n916_), .B2(new_n319_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n319_), .ZN(new_n920_));
  OAI22_X1  g719(.A1(new_n917_), .A2(new_n919_), .B1(new_n920_), .B2(new_n482_), .ZN(new_n921_));
  AOI211_X1 g720(.A(new_n913_), .B(new_n918_), .C1(new_n916_), .C2(new_n319_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n911_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n915_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n865_), .A2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n658_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n918_), .B1(new_n926_), .B2(new_n913_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n917_), .A2(new_n919_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n418_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n927_), .A2(KEYINPUT126), .A3(new_n928_), .A4(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n923_), .A2(new_n930_), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n925_), .B2(new_n636_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n916_), .A2(new_n397_), .A3(new_n746_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1349gat));
  NOR2_X1   g733(.A1(new_n925_), .A2(new_n628_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n935_), .A2(new_n447_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(G183gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n447_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n939_), .B(new_n940_), .C1(G183gat), .C2(new_n935_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n925_), .B2(new_n654_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n916_), .A2(new_n400_), .A3(new_n613_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1351gat));
  NAND3_X1  g744(.A1(new_n894_), .A2(new_n389_), .A3(new_n506_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n658_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n429_), .ZN(G1352gat));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n636_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(new_n430_), .ZN(G1353gat));
  NOR2_X1   g749(.A1(new_n946_), .A2(new_n628_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AND2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n951_), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n954_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  OAI21_X1  g754(.A(G218gat), .B1(new_n946_), .B2(new_n654_), .ZN(new_n956_));
  OR2_X1    g755(.A1(new_n612_), .A2(G218gat), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n946_), .B2(new_n957_), .ZN(G1355gat));
endmodule


