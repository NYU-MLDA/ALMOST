//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_;
  XOR2_X1   g000(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT20), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  INV_X1    g007(.A(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G197gat), .B(G204gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT87), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n215_), .A2(new_n213_), .A3(new_n208_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT23), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n223_), .B(KEYINPUT81), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n225_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT26), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(KEYINPUT26), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n226_), .A2(new_n227_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n228_), .A2(new_n231_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT22), .B(G169gat), .Z(new_n242_));
  OAI211_X1 g041(.A(new_n240_), .B(new_n241_), .C1(G176gat), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n207_), .B1(new_n220_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT19), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n216_), .B(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(new_n218_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n234_), .A2(KEYINPUT80), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(new_n236_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(new_n232_), .C1(KEYINPUT80), .C2(new_n234_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT24), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n229_), .A2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n252_), .A2(new_n222_), .A3(new_n255_), .A4(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n243_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n251_), .A2(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n245_), .A2(new_n248_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n207_), .B1(new_n220_), .B2(new_n259_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n244_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n251_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n248_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n206_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT20), .B1(new_n251_), .B2(new_n264_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n220_), .A2(new_n259_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n247_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n206_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n263_), .A2(new_n248_), .A3(new_n265_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n267_), .A2(new_n273_), .A3(KEYINPUT27), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n263_), .A2(new_n248_), .A3(new_n265_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n248_), .B1(new_n245_), .B2(new_n261_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n206_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT27), .B1(new_n277_), .B2(new_n273_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G85gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G57gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G134gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT83), .ZN(new_n286_));
  XOR2_X1   g085(.A(G113gat), .B(G120gat), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n285_), .A2(KEYINPUT83), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(KEYINPUT83), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n287_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n286_), .A2(KEYINPUT84), .A3(new_n288_), .ZN(new_n295_));
  OR2_X1    g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT85), .ZN(new_n297_));
  XOR2_X1   g096(.A(G155gat), .B(G162gat), .Z(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n296_), .A2(KEYINPUT3), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n296_), .A2(KEYINPUT3), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n298_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n294_), .A2(new_n295_), .B1(new_n303_), .B2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n311_), .A2(KEYINPUT4), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n303_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT4), .B1(new_n311_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G225gat), .A2(G233gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT92), .Z(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n319_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n284_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n284_), .A3(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(KEYINPUT94), .A3(new_n323_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n329_));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT28), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n329_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n220_), .A2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n336_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G22gat), .B(G50gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n333_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n342_), .A3(new_n332_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n294_), .A2(new_n295_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n351_), .A2(new_n352_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n350_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n353_), .A3(new_n349_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n260_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n358_), .A3(new_n259_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT82), .B(G43gat), .Z(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT30), .B(G15gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n362_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n279_), .A2(new_n328_), .A3(new_n348_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n275_), .A2(new_n276_), .A3(new_n206_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n271_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n267_), .A2(new_n273_), .A3(KEYINPUT27), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n326_), .A2(new_n327_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(KEYINPUT95), .A3(new_n348_), .A4(new_n371_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n374_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n345_), .A2(new_n347_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n378_), .A2(new_n327_), .A3(new_n326_), .A4(new_n379_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n371_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n270_), .A2(new_n388_), .A3(new_n272_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n262_), .A2(new_n266_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n324_), .B(new_n389_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n312_), .A2(new_n315_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n283_), .B1(new_n394_), .B2(new_n319_), .ZN(new_n395_));
  OR3_X1    g194(.A1(new_n311_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n321_), .A2(KEYINPUT33), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n277_), .A2(new_n273_), .A3(KEYINPUT91), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n321_), .A2(KEYINPUT33), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT93), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n348_), .B(new_n391_), .C1(new_n399_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n387_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n384_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT71), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT12), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT66), .B(KEYINPUT9), .ZN(new_n407_));
  INV_X1    g206(.A(G92gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT67), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G92gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT9), .ZN(new_n413_));
  OAI21_X1  g212(.A(G85gat), .B1(new_n413_), .B2(new_n408_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n407_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(G85gat), .B2(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G106gat), .ZN(new_n418_));
  INV_X1    g217(.A(G99gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT10), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT10), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT68), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n433_));
  NAND3_X1  g232(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n417_), .A2(new_n426_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n419_), .A3(new_n418_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G85gat), .B(G92gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n432_), .A3(new_n441_), .A4(new_n434_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n444_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n446_), .A2(KEYINPUT8), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n437_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G71gat), .B(G78gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(G57gat), .B(G64gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(KEYINPUT11), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(KEYINPUT11), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n451_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n406_), .B1(new_n457_), .B2(KEYINPUT69), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n459_), .B(KEYINPUT12), .C1(new_n450_), .C2(new_n456_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G230gat), .A2(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT64), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n415_), .A2(new_n416_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n448_), .B1(new_n465_), .B2(new_n426_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n445_), .A3(new_n455_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n457_), .A2(new_n467_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G176gat), .B(G204gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G120gat), .B(G148gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n475_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT13), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT13), .B1(new_n476_), .B2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n405_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n477_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT13), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT71), .A3(new_n478_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G1gat), .A2(G8gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT77), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT14), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n489_), .B2(KEYINPUT14), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G8gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G29gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n498_), .B(KEYINPUT15), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n495_), .B(new_n499_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT79), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n487_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n404_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n501_), .A2(new_n450_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT73), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(KEYINPUT35), .A3(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n499_), .B2(new_n450_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n526_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  INV_X1    g330(.A(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT74), .B(G190gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(KEYINPUT36), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n535_), .B(KEYINPUT36), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n530_), .B2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT37), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n537_), .A2(KEYINPUT75), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n538_), .B(KEYINPUT76), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n530_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n530_), .B2(new_n536_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n543_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n542_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n495_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n456_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G127gat), .B(G155gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT16), .B(G183gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT17), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n557_), .B(KEYINPUT17), .Z(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(new_n553_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT78), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n550_), .A2(new_n563_), .ZN(new_n564_));
  NOR4_X1   g363(.A1(new_n519_), .A2(G1gat), .A3(new_n328_), .A4(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT38), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n486_), .A2(new_n516_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n374_), .A2(new_n383_), .B1(new_n402_), .B2(new_n387_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n540_), .B(KEYINPUT97), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n570_), .A2(new_n562_), .A3(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n573_), .A3(new_n381_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(G1gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n566_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT98), .ZN(G1324gat));
  XNOR2_X1  g376(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(new_n573_), .A3(new_n380_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(G8gat), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT39), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(KEYINPUT39), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n519_), .A2(new_n564_), .ZN(new_n584_));
  INV_X1    g383(.A(G8gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n380_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n578_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n586_), .B(new_n578_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n587_), .A2(new_n589_), .ZN(G1325gat));
  NAND3_X1  g389(.A1(new_n569_), .A2(new_n573_), .A3(new_n371_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(G15gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n591_), .B2(G15gat), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT100), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n593_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT41), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n584_), .A2(new_n603_), .A3(new_n371_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(new_n599_), .A3(KEYINPUT41), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n604_), .A3(new_n605_), .ZN(G1326gat));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n584_), .A2(new_n607_), .A3(new_n385_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n569_), .A2(new_n573_), .A3(new_n385_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G22gat), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT42), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT42), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(G1327gat));
  OR3_X1    g412(.A1(new_n543_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n541_), .B1(new_n614_), .B2(KEYINPUT37), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT43), .B1(new_n550_), .B2(KEYINPUT102), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n404_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n570_), .B2(new_n550_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n569_), .A3(new_n562_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n622_), .A2(new_n569_), .A3(new_n562_), .A4(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n381_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G29gat), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n519_), .A2(new_n563_), .A3(new_n571_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n328_), .A2(G29gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n629_), .B1(new_n631_), .B2(new_n632_), .ZN(G1328gat));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n571_), .A2(new_n563_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n404_), .A2(new_n518_), .A3(new_n634_), .A4(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n279_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT45), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n625_), .A2(new_n380_), .A3(new_n627_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(G36gat), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT104), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n640_), .B(new_n642_), .ZN(G1329gat));
  NAND3_X1  g442(.A1(new_n625_), .A2(new_n371_), .A3(new_n627_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G43gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n371_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n631_), .A2(G43gat), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT47), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(KEYINPUT47), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1330gat));
  NAND3_X1  g451(.A1(new_n625_), .A2(new_n385_), .A3(new_n627_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT105), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n625_), .A2(new_n655_), .A3(new_n385_), .A4(new_n627_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(G50gat), .A3(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n348_), .A2(G50gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n631_), .B2(new_n658_), .ZN(G1331gat));
  NOR2_X1   g458(.A1(new_n570_), .A2(new_n516_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT106), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n487_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n564_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n381_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n486_), .A2(new_n516_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n573_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(G57gat), .A3(new_n381_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n664_), .A2(new_n670_), .A3(new_n671_), .ZN(G1332gat));
  INV_X1    g471(.A(new_n663_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n279_), .A2(G64gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(G64gat), .B1(new_n666_), .B2(new_n279_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT48), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT48), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n673_), .A2(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(G1333gat));
  OR2_X1    g477(.A1(new_n646_), .A2(G71gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(G71gat), .B1(new_n666_), .B2(new_n646_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT49), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT49), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n673_), .A2(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(G1334gat));
  NAND2_X1  g482(.A1(new_n667_), .A2(new_n385_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G78gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT108), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(G78gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT50), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(KEYINPUT50), .A3(new_n688_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n348_), .A2(G78gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n663_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n691_), .B(new_n692_), .C1(new_n694_), .C2(new_n696_), .ZN(G1335gat));
  NAND3_X1  g496(.A1(new_n661_), .A2(new_n487_), .A3(new_n635_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G85gat), .B1(new_n699_), .B2(new_n381_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n481_), .A2(new_n485_), .A3(new_n517_), .A4(new_n562_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n617_), .B2(new_n621_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(new_n381_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n700_), .B1(G85gat), .B2(new_n705_), .ZN(G1336gat));
  AOI21_X1  g505(.A(G92gat), .B1(new_n699_), .B2(new_n380_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n279_), .A2(new_n412_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT111), .Z(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n704_), .B2(new_n709_), .ZN(G1337gat));
  AOI21_X1  g509(.A(new_n419_), .B1(new_n704_), .B2(new_n371_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n424_), .A2(new_n425_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n646_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n699_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT51), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(G1338gat));
  XNOR2_X1  g515(.A(new_n701_), .B(KEYINPUT110), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n616_), .B1(new_n404_), .B2(new_n615_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n570_), .A2(new_n550_), .A3(new_n620_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n385_), .B(new_n717_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G106gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(KEYINPUT113), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n418_), .B1(new_n704_), .B2(new_n385_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n723_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n721_), .A2(KEYINPUT113), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n722_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n698_), .A2(G106gat), .A3(new_n348_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT53), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n721_), .B2(KEYINPUT113), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n725_), .B(new_n723_), .C1(new_n720_), .C2(G106gat), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n732_), .A2(new_n733_), .B1(KEYINPUT113), .B2(new_n721_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  INV_X1    g534(.A(new_n730_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n731_), .A2(new_n737_), .ZN(G1339gat));
  NAND2_X1  g537(.A1(new_n476_), .A2(new_n516_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n464_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT114), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n468_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n455_), .B1(new_n466_), .B2(new_n445_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT12), .B1(new_n744_), .B2(new_n459_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n457_), .A2(KEYINPUT69), .A3(new_n406_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n467_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n463_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(KEYINPUT55), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n742_), .A2(new_n743_), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n748_), .B2(KEYINPUT55), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT114), .B(new_n741_), .C1(new_n747_), .C2(new_n463_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n468_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n754_), .A3(new_n475_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n751_), .A2(new_n754_), .A3(KEYINPUT56), .A4(new_n475_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n739_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n502_), .A2(new_n506_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n505_), .A2(new_n503_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n513_), .A3(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT115), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT115), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n515_), .A3(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n482_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n571_), .B1(new_n759_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n571_), .B(KEYINPUT57), .C1(new_n759_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n476_), .A2(new_n765_), .ZN(new_n772_));
  AND4_X1   g571(.A1(KEYINPUT56), .A2(new_n751_), .A3(new_n754_), .A4(new_n475_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(KEYINPUT116), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n757_), .A2(new_n775_), .A3(new_n758_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n774_), .A2(KEYINPUT58), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT58), .B1(new_n774_), .B2(new_n776_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n550_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n562_), .B1(new_n771_), .B2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n479_), .A2(new_n480_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n550_), .A2(new_n517_), .A3(new_n781_), .A4(new_n563_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT54), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n328_), .A2(new_n380_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n348_), .A3(new_n371_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT117), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(G113gat), .B1(new_n789_), .B2(new_n516_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n517_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n790_), .B1(new_n794_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n486_), .B2(KEYINPUT60), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n796_), .A2(KEYINPUT60), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT118), .ZN(new_n800_));
  OAI21_X1  g599(.A(G120gat), .B1(new_n793_), .B2(new_n486_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1341gat));
  AOI21_X1  g601(.A(G127gat), .B1(new_n789_), .B2(new_n563_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n793_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n563_), .A2(G127gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(G1342gat));
  AOI21_X1  g605(.A(G134gat), .B1(new_n789_), .B2(new_n572_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n615_), .A2(G134gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT119), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n804_), .B2(new_n809_), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n348_), .A2(new_n371_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n785_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n517_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n486_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT120), .B(G148gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n817_), .B(new_n818_), .ZN(G1345gat));
  NOR2_X1   g618(.A1(new_n814_), .A2(new_n562_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT61), .B(G155gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  INV_X1    g621(.A(G162gat), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n814_), .A2(new_n823_), .A3(new_n550_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n813_), .A2(new_n572_), .A3(new_n785_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n823_), .B2(new_n825_), .ZN(G1347gat));
  NOR2_X1   g625(.A1(new_n279_), .A2(new_n381_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n646_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n516_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT121), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n830_), .A2(KEYINPUT121), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n784_), .A2(new_n348_), .A3(new_n831_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT122), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n385_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n831_), .A4(new_n832_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(G169gat), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT62), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n834_), .A2(new_n840_), .A3(G169gat), .A4(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n835_), .A2(new_n829_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n517_), .A2(new_n242_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT123), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1348gat));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n487_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n563_), .ZN(new_n850_));
  MUX2_X1   g649(.A(new_n232_), .B(G183gat), .S(new_n850_), .Z(G1350gat));
  NAND4_X1  g650(.A1(new_n843_), .A2(new_n572_), .A3(new_n236_), .A4(new_n235_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n843_), .A2(new_n615_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n233_), .ZN(G1351gat));
  AOI211_X1 g653(.A(new_n812_), .B(new_n828_), .C1(new_n780_), .C2(new_n783_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n516_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g656(.A1(new_n813_), .A2(new_n487_), .A3(new_n827_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(KEYINPUT124), .A3(new_n487_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(G204gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n858_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT125), .B1(new_n863_), .B2(new_n209_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n860_), .A2(new_n861_), .A3(KEYINPUT125), .A4(G204gat), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1353gat));
  NAND2_X1  g666(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n813_), .A2(new_n563_), .A3(new_n827_), .A4(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT126), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n855_), .A2(new_n871_), .A3(new_n563_), .A4(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1354gat));
  NAND2_X1  g674(.A1(new_n813_), .A2(new_n827_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n532_), .B1(new_n876_), .B2(new_n571_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n855_), .A2(G218gat), .A3(new_n615_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


