//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT23), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n205_), .A2(KEYINPUT77), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT77), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n211_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n214_), .A2(KEYINPUT24), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n209_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(new_n205_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n212_), .B1(new_n224_), .B2(new_n211_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT30), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT30), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(new_n229_), .A3(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G71gat), .B(G99gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G15gat), .B(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n237_), .A2(new_n232_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n232_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n228_), .A2(new_n240_), .A3(new_n230_), .A4(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244_));
  INV_X1    g043(.A(G113gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G120gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT31), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n243_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G141gat), .ZN(new_n250_));
  INV_X1    g049(.A(G148gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(G155gat), .A3(G162gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT80), .Z(new_n256_));
  INV_X1    g055(.A(G155gat), .ZN(new_n257_));
  INV_X1    g056(.A(G162gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(new_n254_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n252_), .B(new_n253_), .C1(new_n256_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT81), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n250_), .B(new_n251_), .C1(new_n263_), .C2(KEYINPUT3), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n265_), .B(KEYINPUT81), .C1(G141gat), .C2(G148gat), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n264_), .A2(new_n266_), .B1(new_n263_), .B2(KEYINPUT3), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n253_), .B(KEYINPUT2), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n260_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n259_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n262_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT29), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT28), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G106gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(KEYINPUT29), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277_));
  INV_X1    g076(.A(G204gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G197gat), .ZN(new_n279_));
  INV_X1    g078(.A(G197gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G204gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n281_), .A3(KEYINPUT83), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n282_), .B(KEYINPUT21), .C1(KEYINPUT83), .C2(new_n281_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n279_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n277_), .B(new_n283_), .C1(new_n286_), .C2(KEYINPUT21), .ZN(new_n287_));
  INV_X1    g086(.A(new_n277_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(KEYINPUT21), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(KEYINPUT82), .A2(G228gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT82), .A2(G228gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(G233gat), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n276_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n294_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n290_), .B(KEYINPUT86), .ZN(new_n299_));
  INV_X1    g098(.A(new_n276_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G22gat), .B(G50gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G78gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n297_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n275_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n274_), .A3(new_n305_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n247_), .A2(new_n271_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n247_), .A2(new_n271_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(KEYINPUT4), .A3(new_n313_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n313_), .A2(KEYINPUT4), .ZN(new_n318_));
  INV_X1    g117(.A(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT0), .B(G57gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G85gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(G1gat), .B(G29gat), .Z(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n316_), .A2(new_n320_), .A3(KEYINPUT33), .A4(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT88), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n325_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT89), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n317_), .A2(new_n318_), .A3(new_n315_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT90), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(KEYINPUT90), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(KEYINPUT89), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .A4(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n316_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  INV_X1    g139(.A(new_n290_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n222_), .A2(new_n215_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n213_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  OAI221_X1 g144(.A(new_n344_), .B1(new_n343_), .B2(new_n225_), .C1(new_n209_), .C2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n341_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT20), .B1(new_n227_), .B2(new_n290_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n340_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n227_), .B2(new_n290_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n341_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n340_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT18), .B(G64gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G92gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  AND3_X1   g157(.A1(new_n349_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n328_), .A2(new_n335_), .A3(new_n338_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n316_), .A2(new_n320_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n324_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n336_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(KEYINPUT91), .A3(new_n324_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n358_), .A2(KEYINPUT32), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n349_), .A2(new_n368_), .A3(new_n354_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n299_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n353_), .B1(new_n370_), .B2(new_n351_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n347_), .A2(new_n348_), .A3(new_n340_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT32), .B(new_n358_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .A4(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n311_), .B1(new_n362_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT92), .B(new_n376_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n358_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n359_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(KEYINPUT27), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n366_), .A2(new_n367_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n310_), .A3(new_n308_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n249_), .B1(new_n375_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n249_), .B1(new_n367_), .B2(new_n366_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n308_), .A2(new_n310_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n381_), .A4(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT93), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n383_), .A2(new_n384_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(KEYINPUT27), .A2(new_n395_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n392_), .A4(new_n391_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT71), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G85gat), .A2(G92gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT66), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT9), .ZN(new_n405_));
  INV_X1    g204(.A(G85gat), .ZN(new_n406_));
  INV_X1    g205(.A(G92gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT9), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n403_), .A3(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT10), .B(G99gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT65), .B(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G99gat), .A2(G106gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n411_), .A2(new_n414_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT7), .ZN(new_n420_));
  INV_X1    g219(.A(G99gat), .ZN(new_n421_));
  INV_X1    g220(.A(G106gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .A4(KEYINPUT67), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT67), .ZN(new_n424_));
  OAI22_X1  g223(.A1(new_n424_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n423_), .A2(new_n425_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT8), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n408_), .A2(new_n428_), .A3(new_n402_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n419_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G50gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G43gat), .ZN(new_n434_));
  INV_X1    g233(.A(G43gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G50gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G36gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G29gat), .ZN(new_n439_));
  INV_X1    g238(.A(G29gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G36gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n434_), .A2(new_n436_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n432_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT15), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT15), .ZN(new_n449_));
  AND4_X1   g248(.A1(new_n434_), .A2(new_n436_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n434_), .A2(new_n436_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n432_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G232gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT34), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n456_), .A2(KEYINPUT35), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n454_), .A2(KEYINPUT69), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT69), .B1(new_n454_), .B2(new_n457_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n456_), .A2(KEYINPUT35), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n457_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n447_), .A2(new_n462_), .A3(new_n453_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT70), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G190gat), .B(G218gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G134gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(new_n258_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT36), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n401_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT71), .B(new_n469_), .C1(new_n460_), .C2(new_n464_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n468_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT36), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(G57gat), .A2(G64gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G57gat), .A2(G64gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G78gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(new_n485_), .A3(new_n480_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n481_), .A2(new_n483_), .A3(KEYINPUT11), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G8gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n202_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G1gat), .A2(G8gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(G15gat), .A2(G22gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G15gat), .A2(G22gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(G1gat), .B2(G8gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n493_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n500_), .A2(new_n497_), .A3(new_n492_), .A4(new_n491_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n489_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT16), .B(G183gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G211gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(G127gat), .B(G155gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  OR3_X1    g309(.A1(new_n505_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(KEYINPUT17), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n478_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n400_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n489_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n432_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n489_), .B(new_n419_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT12), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n432_), .A2(new_n521_), .A3(new_n517_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT64), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n519_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(new_n278_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT5), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n211_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n530_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT13), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n452_), .A2(new_n502_), .A3(new_n448_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n445_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n446_), .A2(new_n502_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n543_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT74), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT74), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n210_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n280_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT75), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n545_), .A2(new_n548_), .A3(KEYINPUT75), .A4(new_n552_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n552_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT76), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT76), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n562_), .B(new_n558_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n538_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n516_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n387_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n202_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT95), .Z(new_n571_));
  NAND3_X1  g370(.A1(new_n475_), .A2(KEYINPUT72), .A3(new_n472_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n401_), .B1(KEYINPUT72), .B2(KEYINPUT37), .ZN(new_n575_));
  INV_X1    g374(.A(new_n465_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n469_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n475_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n514_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n537_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT73), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT73), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n582_), .A2(new_n400_), .A3(new_n565_), .A4(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n202_), .A3(new_n569_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT38), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n571_), .A2(new_n587_), .ZN(G1324gat));
  NAND4_X1  g387(.A1(new_n400_), .A2(new_n567_), .A3(new_n515_), .A4(new_n386_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(KEYINPUT96), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(KEYINPUT96), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(G8gat), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT39), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n590_), .A2(new_n594_), .A3(G8gat), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n585_), .A2(new_n490_), .A3(new_n386_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(KEYINPUT40), .A3(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1325gat));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n249_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n568_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n585_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  INV_X1    g407(.A(G22gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n568_), .B2(new_n311_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT42), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n585_), .A2(new_n609_), .A3(new_n311_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1327gat));
  AOI21_X1  g412(.A(new_n476_), .B1(new_n390_), .B2(new_n399_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n514_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n538_), .A2(new_n566_), .A3(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n440_), .A3(new_n569_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n616_), .B(KEYINPUT97), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n400_), .A2(new_n579_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n572_), .A2(new_n573_), .B1(new_n577_), .B2(new_n475_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n621_), .B2(KEYINPUT98), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n400_), .A2(new_n579_), .A3(new_n622_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n619_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n619_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT99), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n621_), .B(new_n623_), .C1(new_n390_), .C2(new_n399_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n622_), .B1(new_n400_), .B2(new_n579_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n629_), .B(new_n631_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n569_), .A3(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n635_), .A2(KEYINPUT100), .A3(G29gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT100), .B1(new_n635_), .B2(G29gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n618_), .B1(new_n636_), .B2(new_n637_), .ZN(G1328gat));
  OAI211_X1 g437(.A(new_n634_), .B(new_n386_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n617_), .A2(new_n438_), .A3(new_n386_), .A4(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n617_), .A2(new_n438_), .A3(new_n386_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n640_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n639_), .A2(G36gat), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT46), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT102), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT102), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  OAI211_X1 g450(.A(new_n634_), .B(new_n604_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G43gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n617_), .A2(new_n435_), .A3(new_n604_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n655_), .B(new_n657_), .ZN(G1330gat));
  AND4_X1   g457(.A1(G50gat), .A2(new_n628_), .A3(new_n311_), .A4(new_n634_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G50gat), .B1(new_n617_), .B2(new_n311_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g460(.A1(new_n537_), .A2(new_n565_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n400_), .A2(new_n580_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n569_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT104), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n516_), .A2(new_n662_), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT105), .B(G57gat), .Z(new_n667_));
  NOR2_X1   g466(.A1(new_n387_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n665_), .B1(new_n666_), .B2(new_n668_), .ZN(G1332gat));
  INV_X1    g468(.A(G64gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n666_), .B2(new_n386_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT48), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n670_), .A3(new_n386_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1333gat));
  INV_X1    g473(.A(G71gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n666_), .B2(new_n604_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n677_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT49), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n663_), .A2(new_n675_), .A3(new_n604_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(KEYINPUT49), .A3(new_n679_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(G1334gat));
  INV_X1    g484(.A(G78gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n666_), .B2(new_n311_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT50), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n663_), .A2(new_n686_), .A3(new_n311_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1335gat));
  NAND2_X1  g489(.A1(new_n662_), .A2(new_n514_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n614_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT107), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n406_), .A3(new_n569_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT108), .B(new_n692_), .C1(new_n633_), .C2(new_n632_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n387_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n700_), .B2(new_n406_), .ZN(G1336gat));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n407_), .A3(new_n386_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n396_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n407_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT109), .ZN(G1337gat));
  NAND3_X1  g504(.A1(new_n694_), .A2(new_n412_), .A3(new_n604_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n696_), .A2(new_n249_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n421_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g508(.A1(new_n694_), .A2(new_n413_), .A3(new_n311_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G106gat), .B1(new_n696_), .B2(new_n392_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT52), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(KEYINPUT52), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT53), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT53), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n710_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1339gat));
  NAND3_X1  g517(.A1(new_n566_), .A2(KEYINPUT110), .A3(new_n615_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n565_), .B2(new_n514_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n719_), .A2(new_n621_), .A3(new_n537_), .A4(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT54), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n543_), .A2(new_n541_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n540_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n539_), .A2(new_n541_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(new_n551_), .C1(new_n540_), .C2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n557_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n536_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n528_), .A2(KEYINPUT111), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n523_), .B2(KEYINPUT55), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  INV_X1    g531(.A(new_n730_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n732_), .B(new_n733_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n526_), .A2(new_n732_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n534_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(KEYINPUT112), .A2(KEYINPUT56), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n560_), .A2(new_n563_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n530_), .A2(new_n535_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n523_), .A2(KEYINPUT55), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n733_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n523_), .A2(KEYINPUT55), .A3(new_n730_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n736_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n535_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n738_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n741_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n729_), .B1(new_n739_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(KEYINPUT57), .A3(new_n476_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT115), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n476_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n740_), .B1(new_n737_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n757_));
  INV_X1    g556(.A(new_n755_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n746_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n759_), .A3(new_n728_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n756_), .A2(new_n759_), .A3(KEYINPUT58), .A4(new_n728_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n579_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n749_), .A2(new_n765_), .A3(KEYINPUT57), .A4(new_n476_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n751_), .A2(new_n754_), .A3(new_n764_), .A4(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n514_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(new_n514_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n723_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT59), .ZN(new_n772_));
  NOR4_X1   g571(.A1(new_n386_), .A2(new_n311_), .A3(new_n387_), .A4(new_n249_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n767_), .A2(new_n514_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n723_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT59), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT117), .B(G113gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n565_), .A2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT118), .Z(new_n781_));
  NAND3_X1  g580(.A1(new_n774_), .A2(new_n778_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n245_), .B1(new_n777_), .B2(new_n566_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT119), .ZN(G1340gat));
  NAND2_X1  g584(.A1(new_n774_), .A2(new_n778_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G120gat), .B1(new_n786_), .B2(new_n537_), .ZN(new_n787_));
  INV_X1    g586(.A(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n537_), .B2(KEYINPUT60), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT120), .B1(new_n788_), .B2(KEYINPUT60), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n777_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n787_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT121), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n796_), .A3(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1341gat));
  INV_X1    g597(.A(new_n777_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G127gat), .B1(new_n799_), .B2(new_n615_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n774_), .A2(G127gat), .A3(new_n778_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n615_), .ZN(G1342gat));
  INV_X1    g601(.A(new_n478_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n777_), .A2(G134gat), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n774_), .A2(new_n579_), .A3(new_n778_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G134gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT122), .ZN(G1343gat));
  AOI21_X1  g606(.A(new_n604_), .B1(new_n775_), .B2(new_n723_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(new_n569_), .A3(new_n311_), .A4(new_n396_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n566_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(new_n250_), .ZN(G1344gat));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n537_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(new_n251_), .ZN(G1345gat));
  NOR2_X1   g612(.A1(new_n809_), .A2(new_n514_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT61), .B(G155gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1346gat));
  NOR3_X1   g615(.A1(new_n809_), .A2(new_n258_), .A3(new_n621_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n809_), .A2(new_n803_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n258_), .B2(new_n818_), .ZN(G1347gat));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n820_));
  INV_X1    g619(.A(new_n723_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n775_), .A2(KEYINPUT116), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n767_), .A2(new_n768_), .A3(new_n514_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n386_), .A2(new_n391_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n311_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n820_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n771_), .A2(KEYINPUT124), .A3(new_n826_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n565_), .A3(new_n224_), .A4(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n825_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT123), .A3(new_n565_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n825_), .B2(new_n566_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n771_), .A2(new_n392_), .A3(new_n832_), .A4(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n835_), .A2(new_n836_), .A3(G169gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n835_), .B2(G169gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n837_), .B2(new_n838_), .ZN(G1348gat));
  NAND2_X1  g638(.A1(new_n776_), .A2(new_n392_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT125), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n841_), .A2(G176gat), .A3(new_n538_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n828_), .A2(new_n538_), .A3(new_n829_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n842_), .A2(new_n831_), .B1(new_n211_), .B2(new_n843_), .ZN(G1349gat));
  NAND2_X1  g643(.A1(new_n828_), .A2(new_n829_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n514_), .A3(new_n216_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n841_), .A2(new_n615_), .A3(new_n831_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n203_), .B2(new_n847_), .ZN(G1350gat));
  NAND3_X1  g647(.A1(new_n828_), .A2(new_n579_), .A3(new_n829_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G190gat), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n828_), .A2(new_n478_), .A3(new_n217_), .A4(new_n829_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT126), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n854_), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1351gat));
  NOR2_X1   g655(.A1(new_n396_), .A2(new_n388_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n808_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n565_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n280_), .A2(KEYINPUT127), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n280_), .A2(KEYINPUT127), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n862_), .ZN(G1352gat));
  NOR2_X1   g663(.A1(new_n858_), .A2(new_n537_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n278_), .ZN(G1353gat));
  NAND2_X1  g665(.A1(new_n859_), .A2(new_n615_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n868_));
  AND2_X1   g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n867_), .B2(new_n868_), .ZN(G1354gat));
  NOR2_X1   g670(.A1(new_n858_), .A2(new_n803_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n859_), .A2(new_n579_), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n872_), .B(new_n873_), .S(G218gat), .Z(G1355gat));
endmodule


