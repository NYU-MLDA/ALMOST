//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT24), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(KEYINPUT83), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT82), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n209_), .B(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n207_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT79), .B(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT26), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OR3_X1    g021(.A1(new_n222_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT80), .B1(new_n222_), .B2(KEYINPUT26), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n211_), .A2(new_n215_), .A3(new_n219_), .A4(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n203_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n229_));
  AOI21_X1  g028(.A(G176gat), .B1(new_n229_), .B2(G169gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n213_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT85), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n210_), .B2(new_n232_), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n220_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n231_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n227_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n238_), .B(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n246_), .A2(KEYINPUT86), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(KEYINPUT86), .ZN(new_n248_));
  XOR2_X1   g047(.A(G127gat), .B(G134gat), .Z(new_n249_));
  XOR2_X1   g048(.A(G113gat), .B(G120gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT31), .Z(new_n252_));
  OR3_X1    g051(.A1(new_n247_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(KEYINPUT86), .A3(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT88), .B(KEYINPUT3), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT89), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n264_), .A2(KEYINPUT88), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(KEYINPUT88), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n262_), .B(new_n263_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT2), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(G141gat), .A3(G148gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n269_), .A2(new_n271_), .B1(new_n260_), .B2(KEYINPUT3), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n261_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G155gat), .ZN(new_n274_));
  INV_X1    g073(.A(G162gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT87), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(G155gat), .B2(G162gat), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n280_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n260_), .A2(new_n268_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n273_), .A2(new_n281_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT96), .B1(new_n286_), .B2(new_n251_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n273_), .A2(new_n281_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n285_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n288_), .A2(new_n251_), .A3(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n292_), .A3(new_n251_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n256_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n288_), .A2(new_n289_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n251_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n286_), .A2(new_n251_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT96), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n296_), .B1(new_n301_), .B2(new_n293_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n256_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n295_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n295_), .B(new_n313_), .C1(new_n302_), .C2(new_n305_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(KEYINPUT101), .A3(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT4), .B1(new_n291_), .B2(new_n294_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(new_n304_), .A3(new_n303_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT101), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n295_), .A4(new_n313_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n255_), .A2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT28), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G228gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  INV_X1    g128(.A(G204gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT21), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n329_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(G204gat), .A3(new_n335_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT93), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT93), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n334_), .A2(new_n343_), .A3(G204gat), .A4(new_n335_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT92), .B1(new_n329_), .B2(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n330_), .A3(G197gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .A4(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT94), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n344_), .A2(new_n348_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n352_), .A2(KEYINPUT94), .A3(new_n342_), .A4(new_n341_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n339_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n341_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n338_), .A2(new_n342_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n328_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n351_), .A2(new_n353_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n339_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n357_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n360_), .A3(new_n327_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n367_), .A3(KEYINPUT90), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n324_), .A2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n323_), .A2(KEYINPUT90), .A3(new_n362_), .A4(new_n367_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT19), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n213_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT22), .B(G169gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n204_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT26), .B(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n224_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n206_), .A4(new_n212_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT95), .ZN(new_n392_));
  NOR3_X1   g191(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n234_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n387_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n359_), .B2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n238_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n381_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n359_), .B2(new_n395_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n381_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n238_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n379_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n379_), .A3(new_n403_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT27), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(KEYINPUT27), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n391_), .A2(KEYINPUT95), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n394_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n386_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n365_), .A2(new_n357_), .A3(new_n227_), .A4(new_n237_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT20), .A4(new_n401_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n402_), .B(KEYINPUT20), .C1(new_n366_), .C2(new_n415_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n418_), .A2(KEYINPUT100), .B1(new_n419_), .B2(new_n381_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n399_), .B1(new_n366_), .B2(new_n415_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT100), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n401_), .A4(new_n417_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n379_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n410_), .B1(new_n424_), .B2(KEYINPUT103), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n418_), .A2(KEYINPUT100), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n381_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n379_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT103), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n375_), .B(new_n408_), .C1(new_n425_), .C2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT104), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT104), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n409_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n424_), .A2(KEYINPUT103), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n407_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n438_), .B2(new_n375_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n321_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n369_), .A2(new_n370_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n371_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n444_), .A2(new_n372_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n441_), .A2(new_n445_), .A3(new_n408_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT102), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n428_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n398_), .A2(new_n403_), .A3(new_n448_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n320_), .A2(new_n447_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n315_), .A2(new_n450_), .A3(new_n319_), .A4(new_n451_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT102), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n317_), .A2(KEYINPUT33), .A3(new_n295_), .A4(new_n313_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n304_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n303_), .A2(new_n256_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n456_), .B(new_n311_), .C1(new_n302_), .C2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n405_), .A2(new_n455_), .A3(new_n406_), .A4(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n314_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT98), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n314_), .A2(new_n463_), .A3(new_n460_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT99), .B1(new_n459_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n458_), .B1(new_n314_), .B2(new_n460_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n398_), .A2(new_n379_), .A3(new_n403_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n404_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT99), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n452_), .A2(new_n454_), .A3(new_n466_), .A4(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n446_), .B1(new_n472_), .B2(new_n375_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n255_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n440_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G8gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT76), .ZN(new_n477_));
  INV_X1    g276(.A(G22gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n243_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G15gat), .A2(G22gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G1gat), .A2(G8gat), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n479_), .A2(new_n480_), .B1(KEYINPUT14), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n477_), .B(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G29gat), .B(G36gat), .Z(new_n484_));
  XOR2_X1   g283(.A(G43gat), .B(G50gat), .Z(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n483_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n486_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n483_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n483_), .A2(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n489_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT78), .ZN(new_n499_));
  XOR2_X1   g298(.A(G113gat), .B(G141gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT77), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n499_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT6), .ZN(new_n507_));
  OR3_X1    g306(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT66), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n507_), .A2(new_n508_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT8), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT8), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT64), .B(G92gat), .ZN(new_n521_));
  INV_X1    g320(.A(G85gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT9), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n525_));
  INV_X1    g324(.A(G106gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n514_), .A2(KEYINPUT9), .A3(new_n515_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n507_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT65), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n524_), .A2(new_n507_), .A3(new_n530_), .A4(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n518_), .A2(new_n520_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n486_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n493_), .B2(new_n536_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n539_), .A2(new_n540_), .B1(KEYINPUT36), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT72), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n540_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n539_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n538_), .A2(KEYINPUT73), .A3(new_n549_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n544_), .A2(new_n552_), .A3(new_n557_), .A4(new_n553_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT75), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n558_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n562_), .A2(new_n563_), .A3(KEYINPUT37), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n562_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT74), .B1(new_n562_), .B2(KEYINPUT37), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n561_), .A2(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT67), .ZN(new_n569_));
  INV_X1    g368(.A(G64gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G57gat), .ZN(new_n571_));
  INV_X1    g370(.A(G57gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(G64gat), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n573_), .A3(new_n569_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT11), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n576_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT11), .B1(new_n579_), .B2(new_n574_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G71gat), .B(G78gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT11), .B(new_n581_), .C1(new_n579_), .C2(new_n574_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n483_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n588_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n588_), .A2(new_n594_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n568_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n520_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n519_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n532_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n601_), .A2(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n585_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT12), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n518_), .A2(new_n520_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n533_), .A2(new_n535_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n585_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(KEYINPUT68), .A3(KEYINPUT12), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n605_), .A2(KEYINPUT12), .A3(new_n606_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT68), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n609_), .A2(new_n610_), .A3(new_n614_), .A4(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n610_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G120gat), .B(G148gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n620_), .A3(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT70), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(KEYINPUT70), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n618_), .A2(new_n620_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n625_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n629_), .A2(KEYINPUT13), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT13), .B1(new_n629_), .B2(new_n632_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AND4_X1   g434(.A1(new_n475_), .A2(new_n505_), .A3(new_n600_), .A4(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G1gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n320_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n475_), .A2(new_n562_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n505_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n641_), .A2(new_n599_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n637_), .B1(new_n643_), .B2(new_n320_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n639_), .B2(new_n638_), .ZN(G1324gat));
  INV_X1    g445(.A(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n438_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(KEYINPUT105), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(KEYINPUT39), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n438_), .A2(G8gat), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n650_), .A2(new_n654_), .B1(new_n636_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  AOI21_X1  g458(.A(new_n243_), .B1(new_n643_), .B2(new_n474_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n636_), .A2(new_n243_), .A3(new_n474_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(new_n375_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n478_), .B1(new_n643_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n636_), .A2(new_n478_), .A3(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  NAND2_X1  g467(.A1(new_n559_), .A2(new_n599_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT108), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(new_n635_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n475_), .A2(new_n671_), .A3(new_n505_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n475_), .A2(new_n671_), .A3(new_n674_), .A4(new_n505_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n320_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n472_), .A2(new_n375_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n446_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n474_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n320_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n474_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n439_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n438_), .A2(new_n435_), .A3(new_n375_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n678_), .B(new_n568_), .C1(new_n681_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n475_), .A2(KEYINPUT106), .A3(new_n678_), .A4(new_n568_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n475_), .A2(new_n568_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n642_), .A2(new_n598_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n694_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n693_), .A2(KEYINPUT107), .A3(new_n694_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n320_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n677_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  XNOR2_X1  g502(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n697_), .A2(new_n698_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n700_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n695_), .A2(new_n648_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n706_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n438_), .A2(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n673_), .A2(new_n675_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT110), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n673_), .A2(new_n716_), .A3(new_n675_), .A4(new_n713_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(KEYINPUT45), .A3(new_n717_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n705_), .B1(new_n712_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n720_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n718_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n710_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n724_), .B(new_n704_), .C1(new_n725_), .C2(new_n706_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n722_), .A2(new_n726_), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n701_), .A2(G43gat), .A3(new_n474_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  AOI21_X1  g528(.A(G43gat), .B1(new_n676_), .B2(new_n474_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n474_), .A2(G43gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n733_), .B(new_n696_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT47), .B1(new_n734_), .B2(new_n730_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n676_), .B2(new_n664_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n664_), .A2(G50gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n701_), .B2(new_n738_), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n635_), .A2(new_n505_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n598_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n641_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n682_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n475_), .A2(new_n740_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n600_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n572_), .A3(new_n320_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT112), .ZN(G1332gat));
  AOI21_X1  g548(.A(new_n570_), .B1(new_n742_), .B2(new_n648_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT48), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n746_), .A2(new_n570_), .A3(new_n648_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n742_), .B2(new_n474_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n754_), .A3(new_n474_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1334gat));
  INV_X1    g558(.A(G78gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n742_), .B2(new_n664_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT50), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n746_), .A2(new_n760_), .A3(new_n664_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1335gat));
  NAND2_X1  g563(.A1(new_n745_), .A2(new_n670_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT114), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n522_), .A3(new_n320_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n740_), .A2(new_n599_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT115), .Z(new_n769_));
  AND2_X1   g568(.A1(new_n693_), .A2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n320_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n771_), .B2(new_n522_), .ZN(G1336gat));
  AOI21_X1  g571(.A(G92gat), .B1(new_n766_), .B2(new_n648_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n648_), .A2(new_n521_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n770_), .B2(new_n774_), .ZN(G1337gat));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n474_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n474_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(G99gat), .B1(new_n766_), .B2(new_n777_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g578(.A1(new_n766_), .A2(new_n526_), .A3(new_n664_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n693_), .A2(new_n769_), .A3(new_n664_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(G106gat), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n785_), .B(new_n786_), .Z(G1339gat));
  NAND2_X1  g586(.A1(new_n629_), .A2(new_n632_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n503_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n488_), .A2(new_n489_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n495_), .A2(new_n496_), .A3(new_n490_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n498_), .A2(new_n503_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n618_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n536_), .A2(new_n585_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT12), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n536_), .B2(new_n585_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n617_), .A2(new_n614_), .A3(new_n797_), .A4(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n619_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n796_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n618_), .A2(new_n804_), .A3(new_n795_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n618_), .A2(new_n795_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .A4(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n631_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n800_), .A2(new_n619_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n795_), .B2(new_n618_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n618_), .B2(new_n795_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n803_), .B1(new_n813_), .B2(new_n805_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n809_), .C2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n504_), .B1(new_n628_), .B2(new_n627_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n796_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n807_), .A2(new_n818_), .A3(new_n805_), .A4(new_n810_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT119), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n631_), .A3(new_n808_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n821_), .B2(KEYINPUT120), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n794_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n562_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n562_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n814_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n820_), .A2(new_n829_), .A3(new_n631_), .A4(new_n808_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n793_), .A2(new_n792_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(KEYINPUT58), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n567_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n835_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n828_), .A2(new_n837_), .A3(new_n830_), .A4(new_n832_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n827_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n599_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n600_), .A2(new_n504_), .A3(new_n635_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT54), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n434_), .A2(new_n439_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n474_), .A2(new_n320_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n847_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n839_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n836_), .A2(KEYINPUT122), .A3(new_n838_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n826_), .A3(new_n827_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n599_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n852_), .B1(new_n857_), .B2(new_n843_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n851_), .B1(new_n858_), .B2(new_n848_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n504_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n562_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n823_), .B2(new_n562_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n830_), .A2(new_n832_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n805_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n625_), .B1(new_n866_), .B2(new_n803_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n829_), .B1(new_n867_), .B2(new_n820_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n835_), .B1(new_n864_), .B2(new_n868_), .ZN(new_n869_));
  AND4_X1   g668(.A1(KEYINPUT122), .A2(new_n869_), .A3(new_n568_), .A4(new_n838_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT122), .B1(new_n836_), .B2(new_n838_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n598_), .B1(new_n863_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n842_), .B(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n847_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n504_), .A2(G113gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n860_), .B1(new_n876_), .B2(new_n877_), .ZN(G1340gat));
  OAI21_X1  g677(.A(G120gat), .B1(new_n859_), .B2(new_n635_), .ZN(new_n879_));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n635_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(KEYINPUT60), .B2(new_n880_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n876_), .B2(new_n882_), .ZN(G1341gat));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n849_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n876_), .B2(KEYINPUT59), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(new_n598_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n876_), .A2(G127gat), .A3(new_n599_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G127gat), .B1(new_n859_), .B2(new_n599_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  INV_X1    g690(.A(new_n888_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n893_), .ZN(G1342gat));
  OAI21_X1  g693(.A(G134gat), .B1(new_n859_), .B2(new_n567_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n562_), .A2(G134gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n876_), .B2(new_n896_), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n873_), .A2(new_n875_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n474_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n648_), .A2(new_n682_), .A3(new_n375_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n258_), .A3(new_n505_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G141gat), .B1(new_n901_), .B2(new_n504_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1344gat));
  INV_X1    g704(.A(new_n635_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n259_), .A3(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G148gat), .B1(new_n901_), .B2(new_n635_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1345gat));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  OR3_X1    g709(.A1(new_n901_), .A2(new_n599_), .A3(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n901_), .B2(new_n599_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1346gat));
  NAND2_X1  g712(.A1(new_n902_), .A2(new_n559_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n567_), .A2(new_n275_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT124), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n275_), .B1(new_n902_), .B2(new_n916_), .ZN(G1347gat));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n683_), .A2(new_n438_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n664_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n844_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n505_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n918_), .B1(new_n924_), .B2(G169gat), .ZN(new_n925_));
  AOI211_X1 g724(.A(KEYINPUT62), .B(new_n203_), .C1(new_n923_), .C2(new_n505_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n505_), .A2(new_n384_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT125), .Z(new_n928_));
  OAI22_X1  g727(.A1(new_n925_), .A2(new_n926_), .B1(new_n922_), .B2(new_n928_), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n923_), .B2(new_n906_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n898_), .A2(new_n664_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n920_), .A2(new_n204_), .A3(new_n635_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n598_), .A3(new_n919_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n934_), .A2(new_n235_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n922_), .A2(new_n224_), .A3(new_n599_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n936_), .A2(KEYINPUT126), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(KEYINPUT126), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n935_), .A2(new_n937_), .A3(new_n938_), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n922_), .B2(new_n567_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n559_), .A2(new_n388_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n922_), .B2(new_n941_), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n438_), .A2(new_n320_), .A3(new_n375_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n899_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944_), .B2(new_n505_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n899_), .A2(new_n943_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n946_), .A2(new_n329_), .A3(new_n504_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n944_), .A2(new_n330_), .A3(new_n906_), .ZN(new_n949_));
  OAI21_X1  g748(.A(G204gat), .B1(new_n946_), .B2(new_n635_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1353gat));
  AOI21_X1  g750(.A(new_n599_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT127), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n944_), .A2(new_n952_), .A3(new_n954_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n953_), .B(KEYINPUT127), .ZN(new_n956_));
  INV_X1    g755(.A(new_n952_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n946_), .B2(new_n957_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n955_), .A2(new_n958_), .ZN(G1354gat));
  OR3_X1    g758(.A1(new_n946_), .A2(G218gat), .A3(new_n562_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G218gat), .B1(new_n946_), .B2(new_n567_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1355gat));
endmodule


